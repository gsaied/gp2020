
module biasing_fire6_expand1 (
	output [32-1:0] bias_mem [0:256-1]
);

reg [32-1:0] bias_reg_0 = 32'b11111111111111111111111110111111;
reg [32-1:0] bias_reg_1 = 32'b00000000000000000000000000011111;
reg [32-1:0] bias_reg_2 = 32'b11111111111111111111111111111110;
reg [32-1:0] bias_reg_3 = 32'b00000000000000000000000000010101;
reg [32-1:0] bias_reg_4 = 32'b00000000000000000000000000001011;
reg [32-1:0] bias_reg_5 = 32'b11111111111111111111111111111100;
reg [32-1:0] bias_reg_6 = 32'b00000000000000000000000001001000;
reg [32-1:0] bias_reg_7 = 32'b00000000000000000000000000001010;
reg [32-1:0] bias_reg_8 = 32'b00000000000000000000000001010110;
reg [32-1:0] bias_reg_9 = 32'b00000000000000000000000000000110;
reg [32-1:0] bias_reg_10 = 32'b00000000000000000000000000001111;
reg [32-1:0] bias_reg_11 = 32'b00000000000000000000000000111001;
reg [32-1:0] bias_reg_12 = 32'b00000000000000000000000000000110;
reg [32-1:0] bias_reg_13 = 32'b00000000000000000000000000100110;
reg [32-1:0] bias_reg_14 = 32'b00000000000000000000000010000101;
reg [32-1:0] bias_reg_15 = 32'b00000000000000000000000000111111;
reg [32-1:0] bias_reg_16 = 32'b00000000000000000000000000010101;
reg [32-1:0] bias_reg_17 = 32'b00000000000000000000000000001000;
reg [32-1:0] bias_reg_18 = 32'b00000000000000000000000010011101;
reg [32-1:0] bias_reg_19 = 32'b00000000000000000000000001000111;
reg [32-1:0] bias_reg_20 = 32'b00000000000000000000000000111001;
reg [32-1:0] bias_reg_21 = 32'b00000000000000000000000010010101;
reg [32-1:0] bias_reg_22 = 32'b00000000000000000000000000110011;
reg [32-1:0] bias_reg_23 = 32'b00000000000000000000000000100111;
reg [32-1:0] bias_reg_24 = 32'b00000000000000000000000001110111;
reg [32-1:0] bias_reg_25 = 32'b00000000000000000000000000101001;
reg [32-1:0] bias_reg_26 = 32'b11111111111111111111111111010010;
reg [32-1:0] bias_reg_27 = 32'b00000000000000000000000010010001;
reg [32-1:0] bias_reg_28 = 32'b11111111111111111111111111000000;
reg [32-1:0] bias_reg_29 = 32'b00000000000000000000000000110101;
reg [32-1:0] bias_reg_30 = 32'b00000000000000000000000000101110;
reg [32-1:0] bias_reg_31 = 32'b00000000000000000000000000110110;
reg [32-1:0] bias_reg_32 = 32'b00000000000000000000000000010010;
reg [32-1:0] bias_reg_33 = 32'b00000000000000000000000000010010;
reg [32-1:0] bias_reg_34 = 32'b00000000000000000000000000011010;
reg [32-1:0] bias_reg_35 = 32'b11111111111111111111111111101000;
reg [32-1:0] bias_reg_36 = 32'b00000000000000000000000000010111;
reg [32-1:0] bias_reg_37 = 32'b11111111111111111111111111010101;
reg [32-1:0] bias_reg_38 = 32'b00000000000000000000000000011101;
reg [32-1:0] bias_reg_39 = 32'b11111111111111111111111111111010;
reg [32-1:0] bias_reg_40 = 32'b00000000000000000000000010000100;
reg [32-1:0] bias_reg_41 = 32'b00000000000000000000000000010111;
reg [32-1:0] bias_reg_42 = 32'b00000000000000000000000000101011;
reg [32-1:0] bias_reg_43 = 32'b11111111111111111111111111101011;
reg [32-1:0] bias_reg_44 = 32'b00000000000000000000000000101111;
reg [32-1:0] bias_reg_45 = 32'b00000000000000000000000000100111;
reg [32-1:0] bias_reg_46 = 32'b11111111111111111111111111111001;
reg [32-1:0] bias_reg_47 = 32'b00000000000000000000000001100100;
reg [32-1:0] bias_reg_48 = 32'b00000000000000000000000000011010;
reg [32-1:0] bias_reg_49 = 32'b00000000000000000000000000001101;
reg [32-1:0] bias_reg_50 = 32'b00000000000000000000000000001010;
reg [32-1:0] bias_reg_51 = 32'b00000000000000000000000000010001;
reg [32-1:0] bias_reg_52 = 32'b00000000000000000000000000101110;
reg [32-1:0] bias_reg_53 = 32'b00000000000000000000000001100111;
reg [32-1:0] bias_reg_54 = 32'b00000000000000000000000000000110;
reg [32-1:0] bias_reg_55 = 32'b11111111111111111111111111110010;
reg [32-1:0] bias_reg_56 = 32'b00000000000000000000000000101001;
reg [32-1:0] bias_reg_57 = 32'b00000000000000000000000000001110;
reg [32-1:0] bias_reg_58 = 32'b00000000000000000000000000010000;
reg [32-1:0] bias_reg_59 = 32'b00000000000000000000000000000100;
reg [32-1:0] bias_reg_60 = 32'b11111111111111111111111111101111;
reg [32-1:0] bias_reg_61 = 32'b00000000000000000000000000101001;
reg [32-1:0] bias_reg_62 = 32'b00000000000000000000000000011011;
reg [32-1:0] bias_reg_63 = 32'b00000000000000000000000010010101;
reg [32-1:0] bias_reg_64 = 32'b00000000000000000000000000101010;
reg [32-1:0] bias_reg_65 = 32'b00000000000000000000000000100010;
reg [32-1:0] bias_reg_66 = 32'b00000000000000000000000000110010;
reg [32-1:0] bias_reg_67 = 32'b11111111111111111111111111100010;
reg [32-1:0] bias_reg_68 = 32'b11111111111111111111111111110000;
reg [32-1:0] bias_reg_69 = 32'b00000000000000000000000000011011;
reg [32-1:0] bias_reg_70 = 32'b00000000000000000000000000000010;
reg [32-1:0] bias_reg_71 = 32'b00000000000000000000000000010110;
reg [32-1:0] bias_reg_72 = 32'b00000000000000000000000001000001;
reg [32-1:0] bias_reg_73 = 32'b00000000000000000000000000011101;
reg [32-1:0] bias_reg_74 = 32'b00000000000000000000000000011100;
reg [32-1:0] bias_reg_75 = 32'b11111111111111111111111111100001;
reg [32-1:0] bias_reg_76 = 32'b00000000000000000000000001000111;
reg [32-1:0] bias_reg_77 = 32'b00000000000000000000000000011101;
reg [32-1:0] bias_reg_78 = 32'b00000000000000000000000000011110;
reg [32-1:0] bias_reg_79 = 32'b00000000000000000000000000101100;
reg [32-1:0] bias_reg_80 = 32'b00000000000000000000000001110000;
reg [32-1:0] bias_reg_81 = 32'b00000000000000000000000001110011;
reg [32-1:0] bias_reg_82 = 32'b00000000000000000000000000011110;
reg [32-1:0] bias_reg_83 = 32'b00000000000000000000000001101011;
reg [32-1:0] bias_reg_84 = 32'b00000000000000000000000000100111;
reg [32-1:0] bias_reg_85 = 32'b00000000000000000000000000001110;
reg [32-1:0] bias_reg_86 = 32'b11111111111111111111111111111011;
reg [32-1:0] bias_reg_87 = 32'b00000000000000000000000001101101;
reg [32-1:0] bias_reg_88 = 32'b00000000000000000000000000000000;
reg [32-1:0] bias_reg_89 = 32'b00000000000000000000000000001011;
reg [32-1:0] bias_reg_90 = 32'b00000000000000000000000000000111;
reg [32-1:0] bias_reg_91 = 32'b00000000000000000000000000101111;
reg [32-1:0] bias_reg_92 = 32'b11111111111111111111111111011010;
reg [32-1:0] bias_reg_93 = 32'b00000000000000000000000001011001;
reg [32-1:0] bias_reg_94 = 32'b00000000000000000000000001001000;
reg [32-1:0] bias_reg_95 = 32'b00000000000000000000000001111000;
reg [32-1:0] bias_reg_96 = 32'b00000000000000000000000000101110;
reg [32-1:0] bias_reg_97 = 32'b00000000000000000000000000100001;
reg [32-1:0] bias_reg_98 = 32'b00000000000000000000000010010000;
reg [32-1:0] bias_reg_99 = 32'b00000000000000000000000000000010;
reg [32-1:0] bias_reg_100 = 32'b00000000000000000000000000001011;
reg [32-1:0] bias_reg_101 = 32'b00000000000000000000000010101001;
reg [32-1:0] bias_reg_102 = 32'b00000000000000000000000000001111;
reg [32-1:0] bias_reg_103 = 32'b11111111111111111111111111111111;
reg [32-1:0] bias_reg_104 = 32'b00000000000000000000000000000001;
reg [32-1:0] bias_reg_105 = 32'b00000000000000000000000000011100;
reg [32-1:0] bias_reg_106 = 32'b00000000000000000000000001010000;
reg [32-1:0] bias_reg_107 = 32'b00000000000000000000000000101101;
reg [32-1:0] bias_reg_108 = 32'b00000000000000000000000000111100;
reg [32-1:0] bias_reg_109 = 32'b00000000000000000000000000001111;
reg [32-1:0] bias_reg_110 = 32'b00000000000000000000000001010011;
reg [32-1:0] bias_reg_111 = 32'b00000000000000000000000000110000;
reg [32-1:0] bias_reg_112 = 32'b00000000000000000000000000100011;
reg [32-1:0] bias_reg_113 = 32'b00000000000000000000000000101111;
reg [32-1:0] bias_reg_114 = 32'b11111111111111111111111111110001;
reg [32-1:0] bias_reg_115 = 32'b00000000000000000000000000101010;
reg [32-1:0] bias_reg_116 = 32'b00000000000000000000000000000001;
reg [32-1:0] bias_reg_117 = 32'b00000000000000000000000000111110;
reg [32-1:0] bias_reg_118 = 32'b00000000000000000000000000110111;
reg [32-1:0] bias_reg_119 = 32'b00000000000000000000000000011001;
reg [32-1:0] bias_reg_120 = 32'b00000000000000000000000001011010;
reg [32-1:0] bias_reg_121 = 32'b11111111111111111111111111101111;
reg [32-1:0] bias_reg_122 = 32'b11111111111111111111111111110100;
reg [32-1:0] bias_reg_123 = 32'b00000000000000000000000001000111;
reg [32-1:0] bias_reg_124 = 32'b00000000000000000000000000101101;
reg [32-1:0] bias_reg_125 = 32'b00000000000000000000000001000011;
reg [32-1:0] bias_reg_126 = 32'b00000000000000000000000001001101;
reg [32-1:0] bias_reg_127 = 32'b00000000000000000000000001000011;
reg [32-1:0] bias_reg_128 = 32'b11111111111111111111111101111001;
reg [32-1:0] bias_reg_129 = 32'b00000000000000000000000000010010;
reg [32-1:0] bias_reg_130 = 32'b00000000000000000000000000010011;
reg [32-1:0] bias_reg_131 = 32'b00000000000000000000000000101001;
reg [32-1:0] bias_reg_132 = 32'b00000000000000000000000000011110;
reg [32-1:0] bias_reg_133 = 32'b00000000000000000000000001001000;
reg [32-1:0] bias_reg_134 = 32'b00000000000000000000000000111010;
reg [32-1:0] bias_reg_135 = 32'b00000000000000000000000001100001;
reg [32-1:0] bias_reg_136 = 32'b00000000000000000000000000100101;
reg [32-1:0] bias_reg_137 = 32'b00000000000000000000000000010101;
reg [32-1:0] bias_reg_138 = 32'b11111111111111111111111111101111;
reg [32-1:0] bias_reg_139 = 32'b00000000000000000000000001001010;
reg [32-1:0] bias_reg_140 = 32'b00000000000000000000000100001011;
reg [32-1:0] bias_reg_141 = 32'b00000000000000000000000000000110;
reg [32-1:0] bias_reg_142 = 32'b00000000000000000000000000110010;
reg [32-1:0] bias_reg_143 = 32'b00000000000000000000000000000000;
reg [32-1:0] bias_reg_144 = 32'b00000000000000000000000000000010;
reg [32-1:0] bias_reg_145 = 32'b00000000000000000000000001100111;
reg [32-1:0] bias_reg_146 = 32'b00000000000000000000000000010110;
reg [32-1:0] bias_reg_147 = 32'b00000000000000000000000000111001;
reg [32-1:0] bias_reg_148 = 32'b11111111111111111111111111111101;
reg [32-1:0] bias_reg_149 = 32'b11111111111111111111111110101000;
reg [32-1:0] bias_reg_150 = 32'b00000000000000000000000000111100;
reg [32-1:0] bias_reg_151 = 32'b00000000000000000000000000101100;
reg [32-1:0] bias_reg_152 = 32'b11111111111111111111111111001110;
reg [32-1:0] bias_reg_153 = 32'b00000000000000000000000000010000;
reg [32-1:0] bias_reg_154 = 32'b00000000000000000000000000001001;
reg [32-1:0] bias_reg_155 = 32'b00000000000000000000000000110010;
reg [32-1:0] bias_reg_156 = 32'b00000000000000000000000000000100;
reg [32-1:0] bias_reg_157 = 32'b00000000000000000000000000110000;
reg [32-1:0] bias_reg_158 = 32'b00000000000000000000000000110011;
reg [32-1:0] bias_reg_159 = 32'b00000000000000000000000000000011;
reg [32-1:0] bias_reg_160 = 32'b00000000000000000000000001000010;
reg [32-1:0] bias_reg_161 = 32'b00000000000000000000000000011011;
reg [32-1:0] bias_reg_162 = 32'b00000000000000000000000001111010;
reg [32-1:0] bias_reg_163 = 32'b11111111111111111111111111110100;
reg [32-1:0] bias_reg_164 = 32'b11111111111111111111111111101001;
reg [32-1:0] bias_reg_165 = 32'b11111111111111111111111111111101;
reg [32-1:0] bias_reg_166 = 32'b00000000000000000000000000100010;
reg [32-1:0] bias_reg_167 = 32'b11111111111111111111111111100110;
reg [32-1:0] bias_reg_168 = 32'b11111111111111111111111111110010;
reg [32-1:0] bias_reg_169 = 32'b00000000000000000000000001101101;
reg [32-1:0] bias_reg_170 = 32'b00000000000000000000000001100111;
reg [32-1:0] bias_reg_171 = 32'b00000000000000000000000000111010;
reg [32-1:0] bias_reg_172 = 32'b00000000000000000000000000010101;
reg [32-1:0] bias_reg_173 = 32'b00000000000000000000000001000010;
reg [32-1:0] bias_reg_174 = 32'b11111111111111111111111111110010;
reg [32-1:0] bias_reg_175 = 32'b00000000000000000000000000110100;
reg [32-1:0] bias_reg_176 = 32'b00000000000000000000000001000001;
reg [32-1:0] bias_reg_177 = 32'b00000000000000000000000000110110;
reg [32-1:0] bias_reg_178 = 32'b00000000000000000000000000101010;
reg [32-1:0] bias_reg_179 = 32'b00000000000000000000000001001111;
reg [32-1:0] bias_reg_180 = 32'b00000000000000000000000000100010;
reg [32-1:0] bias_reg_181 = 32'b00000000000000000000000000110001;
reg [32-1:0] bias_reg_182 = 32'b11111111111111111111111111100000;
reg [32-1:0] bias_reg_183 = 32'b00000000000000000000000000000001;
reg [32-1:0] bias_reg_184 = 32'b00000000000000000000000001101111;
reg [32-1:0] bias_reg_185 = 32'b00000000000000000000000000110001;
reg [32-1:0] bias_reg_186 = 32'b00000000000000000000000000010110;
reg [32-1:0] bias_reg_187 = 32'b11111111111111111111111111111101;
reg [32-1:0] bias_reg_188 = 32'b11111111111111111111111111111100;
reg [32-1:0] bias_reg_189 = 32'b00000000000000000000000000010001;
reg [32-1:0] bias_reg_190 = 32'b11111111111111111111111111110101;
reg [32-1:0] bias_reg_191 = 32'b11111111111111111111111111111111;
reg [32-1:0] bias_reg_192 = 32'b00000000000000000000000000100110;
reg [32-1:0] bias_reg_193 = 32'b00000000000000000000000001001101;
reg [32-1:0] bias_reg_194 = 32'b11111111111111111111111111011100;
reg [32-1:0] bias_reg_195 = 32'b00000000000000000000000000010101;
reg [32-1:0] bias_reg_196 = 32'b11111111111111111111111111111001;
reg [32-1:0] bias_reg_197 = 32'b00000000000000000000000000011001;
reg [32-1:0] bias_reg_198 = 32'b00000000000000000000000000000010;
reg [32-1:0] bias_reg_199 = 32'b00000000000000000000000000110011;
reg [32-1:0] bias_reg_200 = 32'b11111111111111111111111111011100;
reg [32-1:0] bias_reg_201 = 32'b11111111111111111111111111001011;
reg [32-1:0] bias_reg_202 = 32'b00000000000000000000000001101011;
reg [32-1:0] bias_reg_203 = 32'b00000000000000000000000001111001;
reg [32-1:0] bias_reg_204 = 32'b00000000000000000000000000010011;
reg [32-1:0] bias_reg_205 = 32'b00000000000000000000000001001001;
reg [32-1:0] bias_reg_206 = 32'b00000000000000000000000001001010;
reg [32-1:0] bias_reg_207 = 32'b00000000000000000000000011100100;
reg [32-1:0] bias_reg_208 = 32'b00000000000000000000000001001010;
reg [32-1:0] bias_reg_209 = 32'b00000000000000000000000001101011;
reg [32-1:0] bias_reg_210 = 32'b00000000000000000000000001000010;
reg [32-1:0] bias_reg_211 = 32'b00000000000000000000000000001000;
reg [32-1:0] bias_reg_212 = 32'b11111111111111111111111111101101;
reg [32-1:0] bias_reg_213 = 32'b00000000000000000000000001011100;
reg [32-1:0] bias_reg_214 = 32'b00000000000000000000000001001111;
reg [32-1:0] bias_reg_215 = 32'b11111111111111111111111111010010;
reg [32-1:0] bias_reg_216 = 32'b00000000000000000000000010001001;
reg [32-1:0] bias_reg_217 = 32'b11111111111111111111111111100110;
reg [32-1:0] bias_reg_218 = 32'b00000000000000000000000000111101;
reg [32-1:0] bias_reg_219 = 32'b00000000000000000000000001010100;
reg [32-1:0] bias_reg_220 = 32'b11111111111111111111111111111000;
reg [32-1:0] bias_reg_221 = 32'b00000000000000000000000000100010;
reg [32-1:0] bias_reg_222 = 32'b00000000000000000000000001010010;
reg [32-1:0] bias_reg_223 = 32'b00000000000000000000000001010101;
reg [32-1:0] bias_reg_224 = 32'b00000000000000000000000000001110;
reg [32-1:0] bias_reg_225 = 32'b00000000000000000000000000010010;
reg [32-1:0] bias_reg_226 = 32'b11111111111111111111111111100101;
reg [32-1:0] bias_reg_227 = 32'b11111111111111111111111111101100;
reg [32-1:0] bias_reg_228 = 32'b11111111111111111111111111011010;
reg [32-1:0] bias_reg_229 = 32'b00000000000000000000000001000101;
reg [32-1:0] bias_reg_230 = 32'b00000000000000000000000000110111;
reg [32-1:0] bias_reg_231 = 32'b00000000000000000000000000011101;
reg [32-1:0] bias_reg_232 = 32'b00000000000000000000000000011010;
reg [32-1:0] bias_reg_233 = 32'b00000000000000000000000000001011;
reg [32-1:0] bias_reg_234 = 32'b00000000000000000000000000011010;
reg [32-1:0] bias_reg_235 = 32'b00000000000000000000000000101000;
reg [32-1:0] bias_reg_236 = 32'b11111111111111111111111111000000;
reg [32-1:0] bias_reg_237 = 32'b00000000000000000000000000001001;
reg [32-1:0] bias_reg_238 = 32'b00000000000000000000000000101010;
reg [32-1:0] bias_reg_239 = 32'b00000000000000000000000001000101;
reg [32-1:0] bias_reg_240 = 32'b00000000000000000000000001100100;
reg [32-1:0] bias_reg_241 = 32'b00000000000000000000000000011100;
reg [32-1:0] bias_reg_242 = 32'b00000000000000000000000001100100;
reg [32-1:0] bias_reg_243 = 32'b11111111111111111111111111011001;
reg [32-1:0] bias_reg_244 = 32'b00000000000000000000000000101000;
reg [32-1:0] bias_reg_245 = 32'b00000000000000000000000000000110;
reg [32-1:0] bias_reg_246 = 32'b11111111111111111111111111111001;
reg [32-1:0] bias_reg_247 = 32'b00000000000000000000000001110010;
reg [32-1:0] bias_reg_248 = 32'b00000000000000000000000000101001;
reg [32-1:0] bias_reg_249 = 32'b00000000000000000000000001001110;
reg [32-1:0] bias_reg_250 = 32'b11111111111111111111111111101011;
reg [32-1:0] bias_reg_251 = 32'b00000000000000000000000001000000;
reg [32-1:0] bias_reg_252 = 32'b00000000000000000000000001000101;
reg [32-1:0] bias_reg_253 = 32'b00000000000000000000000001011010;
reg [32-1:0] bias_reg_254 = 32'b11111111111111111111111111101100;
reg [32-1:0] bias_reg_255 = 32'b00000000000000000000000001111010;
assign bias_mem[0] = bias_reg_0;
assign bias_mem[1] = bias_reg_1;
assign bias_mem[2] = bias_reg_2;
assign bias_mem[3] = bias_reg_3;
assign bias_mem[4] = bias_reg_4;
assign bias_mem[5] = bias_reg_5;
assign bias_mem[6] = bias_reg_6;
assign bias_mem[7] = bias_reg_7;
assign bias_mem[8] = bias_reg_8;
assign bias_mem[9] = bias_reg_9;
assign bias_mem[10] = bias_reg_10;
assign bias_mem[11] = bias_reg_11;
assign bias_mem[12] = bias_reg_12;
assign bias_mem[13] = bias_reg_13;
assign bias_mem[14] = bias_reg_14;
assign bias_mem[15] = bias_reg_15;
assign bias_mem[16] = bias_reg_16;
assign bias_mem[17] = bias_reg_17;
assign bias_mem[18] = bias_reg_18;
assign bias_mem[19] = bias_reg_19;
assign bias_mem[20] = bias_reg_20;
assign bias_mem[21] = bias_reg_21;
assign bias_mem[22] = bias_reg_22;
assign bias_mem[23] = bias_reg_23;
assign bias_mem[24] = bias_reg_24;
assign bias_mem[25] = bias_reg_25;
assign bias_mem[26] = bias_reg_26;
assign bias_mem[27] = bias_reg_27;
assign bias_mem[28] = bias_reg_28;
assign bias_mem[29] = bias_reg_29;
assign bias_mem[30] = bias_reg_30;
assign bias_mem[31] = bias_reg_31;
assign bias_mem[32] = bias_reg_32;
assign bias_mem[33] = bias_reg_33;
assign bias_mem[34] = bias_reg_34;
assign bias_mem[35] = bias_reg_35;
assign bias_mem[36] = bias_reg_36;
assign bias_mem[37] = bias_reg_37;
assign bias_mem[38] = bias_reg_38;
assign bias_mem[39] = bias_reg_39;
assign bias_mem[40] = bias_reg_40;
assign bias_mem[41] = bias_reg_41;
assign bias_mem[42] = bias_reg_42;
assign bias_mem[43] = bias_reg_43;
assign bias_mem[44] = bias_reg_44;
assign bias_mem[45] = bias_reg_45;
assign bias_mem[46] = bias_reg_46;
assign bias_mem[47] = bias_reg_47;
assign bias_mem[48] = bias_reg_48;
assign bias_mem[49] = bias_reg_49;
assign bias_mem[50] = bias_reg_50;
assign bias_mem[51] = bias_reg_51;
assign bias_mem[52] = bias_reg_52;
assign bias_mem[53] = bias_reg_53;
assign bias_mem[54] = bias_reg_54;
assign bias_mem[55] = bias_reg_55;
assign bias_mem[56] = bias_reg_56;
assign bias_mem[57] = bias_reg_57;
assign bias_mem[58] = bias_reg_58;
assign bias_mem[59] = bias_reg_59;
assign bias_mem[60] = bias_reg_60;
assign bias_mem[61] = bias_reg_61;
assign bias_mem[62] = bias_reg_62;
assign bias_mem[63] = bias_reg_63;
assign bias_mem[64] = bias_reg_64;
assign bias_mem[65] = bias_reg_65;
assign bias_mem[66] = bias_reg_66;
assign bias_mem[67] = bias_reg_67;
assign bias_mem[68] = bias_reg_68;
assign bias_mem[69] = bias_reg_69;
assign bias_mem[70] = bias_reg_70;
assign bias_mem[71] = bias_reg_71;
assign bias_mem[72] = bias_reg_72;
assign bias_mem[73] = bias_reg_73;
assign bias_mem[74] = bias_reg_74;
assign bias_mem[75] = bias_reg_75;
assign bias_mem[76] = bias_reg_76;
assign bias_mem[77] = bias_reg_77;
assign bias_mem[78] = bias_reg_78;
assign bias_mem[79] = bias_reg_79;
assign bias_mem[80] = bias_reg_80;
assign bias_mem[81] = bias_reg_81;
assign bias_mem[82] = bias_reg_82;
assign bias_mem[83] = bias_reg_83;
assign bias_mem[84] = bias_reg_84;
assign bias_mem[85] = bias_reg_85;
assign bias_mem[86] = bias_reg_86;
assign bias_mem[87] = bias_reg_87;
assign bias_mem[88] = bias_reg_88;
assign bias_mem[89] = bias_reg_89;
assign bias_mem[90] = bias_reg_90;
assign bias_mem[91] = bias_reg_91;
assign bias_mem[92] = bias_reg_92;
assign bias_mem[93] = bias_reg_93;
assign bias_mem[94] = bias_reg_94;
assign bias_mem[95] = bias_reg_95;
assign bias_mem[96] = bias_reg_96;
assign bias_mem[97] = bias_reg_97;
assign bias_mem[98] = bias_reg_98;
assign bias_mem[99] = bias_reg_99;
assign bias_mem[100] = bias_reg_100;
assign bias_mem[101] = bias_reg_101;
assign bias_mem[102] = bias_reg_102;
assign bias_mem[103] = bias_reg_103;
assign bias_mem[104] = bias_reg_104;
assign bias_mem[105] = bias_reg_105;
assign bias_mem[106] = bias_reg_106;
assign bias_mem[107] = bias_reg_107;
assign bias_mem[108] = bias_reg_108;
assign bias_mem[109] = bias_reg_109;
assign bias_mem[110] = bias_reg_110;
assign bias_mem[111] = bias_reg_111;
assign bias_mem[112] = bias_reg_112;
assign bias_mem[113] = bias_reg_113;
assign bias_mem[114] = bias_reg_114;
assign bias_mem[115] = bias_reg_115;
assign bias_mem[116] = bias_reg_116;
assign bias_mem[117] = bias_reg_117;
assign bias_mem[118] = bias_reg_118;
assign bias_mem[119] = bias_reg_119;
assign bias_mem[120] = bias_reg_120;
assign bias_mem[121] = bias_reg_121;
assign bias_mem[122] = bias_reg_122;
assign bias_mem[123] = bias_reg_123;
assign bias_mem[124] = bias_reg_124;
assign bias_mem[125] = bias_reg_125;
assign bias_mem[126] = bias_reg_126;
assign bias_mem[127] = bias_reg_127;
assign bias_mem[128] = bias_reg_128;
assign bias_mem[129] = bias_reg_129;
assign bias_mem[130] = bias_reg_130;
assign bias_mem[131] = bias_reg_131;
assign bias_mem[132] = bias_reg_132;
assign bias_mem[133] = bias_reg_133;
assign bias_mem[134] = bias_reg_134;
assign bias_mem[135] = bias_reg_135;
assign bias_mem[136] = bias_reg_136;
assign bias_mem[137] = bias_reg_137;
assign bias_mem[138] = bias_reg_138;
assign bias_mem[139] = bias_reg_139;
assign bias_mem[140] = bias_reg_140;
assign bias_mem[141] = bias_reg_141;
assign bias_mem[142] = bias_reg_142;
assign bias_mem[143] = bias_reg_143;
assign bias_mem[144] = bias_reg_144;
assign bias_mem[145] = bias_reg_145;
assign bias_mem[146] = bias_reg_146;
assign bias_mem[147] = bias_reg_147;
assign bias_mem[148] = bias_reg_148;
assign bias_mem[149] = bias_reg_149;
assign bias_mem[150] = bias_reg_150;
assign bias_mem[151] = bias_reg_151;
assign bias_mem[152] = bias_reg_152;
assign bias_mem[153] = bias_reg_153;
assign bias_mem[154] = bias_reg_154;
assign bias_mem[155] = bias_reg_155;
assign bias_mem[156] = bias_reg_156;
assign bias_mem[157] = bias_reg_157;
assign bias_mem[158] = bias_reg_158;
assign bias_mem[159] = bias_reg_159;
assign bias_mem[160] = bias_reg_160;
assign bias_mem[161] = bias_reg_161;
assign bias_mem[162] = bias_reg_162;
assign bias_mem[163] = bias_reg_163;
assign bias_mem[164] = bias_reg_164;
assign bias_mem[165] = bias_reg_165;
assign bias_mem[166] = bias_reg_166;
assign bias_mem[167] = bias_reg_167;
assign bias_mem[168] = bias_reg_168;
assign bias_mem[169] = bias_reg_169;
assign bias_mem[170] = bias_reg_170;
assign bias_mem[171] = bias_reg_171;
assign bias_mem[172] = bias_reg_172;
assign bias_mem[173] = bias_reg_173;
assign bias_mem[174] = bias_reg_174;
assign bias_mem[175] = bias_reg_175;
assign bias_mem[176] = bias_reg_176;
assign bias_mem[177] = bias_reg_177;
assign bias_mem[178] = bias_reg_178;
assign bias_mem[179] = bias_reg_179;
assign bias_mem[180] = bias_reg_180;
assign bias_mem[181] = bias_reg_181;
assign bias_mem[182] = bias_reg_182;
assign bias_mem[183] = bias_reg_183;
assign bias_mem[184] = bias_reg_184;
assign bias_mem[185] = bias_reg_185;
assign bias_mem[186] = bias_reg_186;
assign bias_mem[187] = bias_reg_187;
assign bias_mem[188] = bias_reg_188;
assign bias_mem[189] = bias_reg_189;
assign bias_mem[190] = bias_reg_190;
assign bias_mem[191] = bias_reg_191;
assign bias_mem[192] = bias_reg_192;
assign bias_mem[193] = bias_reg_193;
assign bias_mem[194] = bias_reg_194;
assign bias_mem[195] = bias_reg_195;
assign bias_mem[196] = bias_reg_196;
assign bias_mem[197] = bias_reg_197;
assign bias_mem[198] = bias_reg_198;
assign bias_mem[199] = bias_reg_199;
assign bias_mem[200] = bias_reg_200;
assign bias_mem[201] = bias_reg_201;
assign bias_mem[202] = bias_reg_202;
assign bias_mem[203] = bias_reg_203;
assign bias_mem[204] = bias_reg_204;
assign bias_mem[205] = bias_reg_205;
assign bias_mem[206] = bias_reg_206;
assign bias_mem[207] = bias_reg_207;
assign bias_mem[208] = bias_reg_208;
assign bias_mem[209] = bias_reg_209;
assign bias_mem[210] = bias_reg_210;
assign bias_mem[211] = bias_reg_211;
assign bias_mem[212] = bias_reg_212;
assign bias_mem[213] = bias_reg_213;
assign bias_mem[214] = bias_reg_214;
assign bias_mem[215] = bias_reg_215;
assign bias_mem[216] = bias_reg_216;
assign bias_mem[217] = bias_reg_217;
assign bias_mem[218] = bias_reg_218;
assign bias_mem[219] = bias_reg_219;
assign bias_mem[220] = bias_reg_220;
assign bias_mem[221] = bias_reg_221;
assign bias_mem[222] = bias_reg_222;
assign bias_mem[223] = bias_reg_223;
assign bias_mem[224] = bias_reg_224;
assign bias_mem[225] = bias_reg_225;
assign bias_mem[226] = bias_reg_226;
assign bias_mem[227] = bias_reg_227;
assign bias_mem[228] = bias_reg_228;
assign bias_mem[229] = bias_reg_229;
assign bias_mem[230] = bias_reg_230;
assign bias_mem[231] = bias_reg_231;
assign bias_mem[232] = bias_reg_232;
assign bias_mem[233] = bias_reg_233;
assign bias_mem[234] = bias_reg_234;
assign bias_mem[235] = bias_reg_235;
assign bias_mem[236] = bias_reg_236;
assign bias_mem[237] = bias_reg_237;
assign bias_mem[238] = bias_reg_238;
assign bias_mem[239] = bias_reg_239;
assign bias_mem[240] = bias_reg_240;
assign bias_mem[241] = bias_reg_241;
assign bias_mem[242] = bias_reg_242;
assign bias_mem[243] = bias_reg_243;
assign bias_mem[244] = bias_reg_244;
assign bias_mem[245] = bias_reg_245;
assign bias_mem[246] = bias_reg_246;
assign bias_mem[247] = bias_reg_247;
assign bias_mem[248] = bias_reg_248;
assign bias_mem[249] = bias_reg_249;
assign bias_mem[250] = bias_reg_250;
assign bias_mem[251] = bias_reg_251;
assign bias_mem[252] = bias_reg_252;
assign bias_mem[253] = bias_reg_253;
assign bias_mem[254] = bias_reg_254;
assign bias_mem[255] = bias_reg_255;
endmodule
