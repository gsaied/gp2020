
module biasing_fire7_squeeze (
	output [32-1:0] bias_mem [0:64-1]
);

reg [32-1:0] bias_reg_0 = 32'b11111111111111111111111101000101;
reg [32-1:0] bias_reg_1 = 32'b11111111111111111111111111101100;
reg [32-1:0] bias_reg_2 = 32'b00000000000000000000000000110101;
reg [32-1:0] bias_reg_3 = 32'b00000000000000000000000000101001;
reg [32-1:0] bias_reg_4 = 32'b11111111111111111111111110000110;
reg [32-1:0] bias_reg_5 = 32'b00000000000000000000000001000011;
reg [32-1:0] bias_reg_6 = 32'b00000000000000000000000001001001;
reg [32-1:0] bias_reg_7 = 32'b11111111111111111111111110100000;
reg [32-1:0] bias_reg_8 = 32'b11111111111111111111111110101110;
reg [32-1:0] bias_reg_9 = 32'b11111111111111111111111111001100;
reg [32-1:0] bias_reg_10 = 32'b11111111111111111111111101011000;
reg [32-1:0] bias_reg_11 = 32'b11111111111111111111111011110010;
reg [32-1:0] bias_reg_12 = 32'b00000000000000000000000001011101;
reg [32-1:0] bias_reg_13 = 32'b11111111111111111111111111010111;
reg [32-1:0] bias_reg_14 = 32'b11111111111111111111111011111011;
reg [32-1:0] bias_reg_15 = 32'b00000000000000000000000001101001;
reg [32-1:0] bias_reg_16 = 32'b00000000000000000000000001101000;
reg [32-1:0] bias_reg_17 = 32'b11111111111111111111111101101001;
reg [32-1:0] bias_reg_18 = 32'b00000000000000000000000100101111;
reg [32-1:0] bias_reg_19 = 32'b00000000000000000000000001010000;
reg [32-1:0] bias_reg_20 = 32'b11111111111111111111111110001010;
reg [32-1:0] bias_reg_21 = 32'b00000000000000000000000000010111;
reg [32-1:0] bias_reg_22 = 32'b00000000000000000000000001011111;
reg [32-1:0] bias_reg_23 = 32'b00000000000000000000000011001000;
reg [32-1:0] bias_reg_24 = 32'b11111111111111111111111110100001;
reg [32-1:0] bias_reg_25 = 32'b11111111111111111111111101111101;
reg [32-1:0] bias_reg_26 = 32'b00000000000000000000000100110101;
reg [32-1:0] bias_reg_27 = 32'b00000000000000000000000001011000;
reg [32-1:0] bias_reg_28 = 32'b00000000000000000000000010111000;
reg [32-1:0] bias_reg_29 = 32'b00000000000000000000000001011100;
reg [32-1:0] bias_reg_30 = 32'b00000000000000000000000010000110;
reg [32-1:0] bias_reg_31 = 32'b11111111111111111111111111010101;
reg [32-1:0] bias_reg_32 = 32'b00000000000000000000000011001111;
reg [32-1:0] bias_reg_33 = 32'b00000000000000000000000000000011;
reg [32-1:0] bias_reg_34 = 32'b11111111111111111111111110111000;
reg [32-1:0] bias_reg_35 = 32'b00000000000000000000000011000111;
reg [32-1:0] bias_reg_36 = 32'b11111111111111111111110000000111;
reg [32-1:0] bias_reg_37 = 32'b00000000000000000000010101001101;
reg [32-1:0] bias_reg_38 = 32'b00000000000000000000000001100101;
reg [32-1:0] bias_reg_39 = 32'b00000000000000000000000000101001;
reg [32-1:0] bias_reg_40 = 32'b00000000000000000000000001000110;
reg [32-1:0] bias_reg_41 = 32'b00000000000000000000000000110111;
reg [32-1:0] bias_reg_42 = 32'b11111111111111111111111111100000;
reg [32-1:0] bias_reg_43 = 32'b00000000000000000000000000100100;
reg [32-1:0] bias_reg_44 = 32'b00000000000000000000000001010100;
reg [32-1:0] bias_reg_45 = 32'b11111111111111111111111111101101;
reg [32-1:0] bias_reg_46 = 32'b00000000000000000000000000001011;
reg [32-1:0] bias_reg_47 = 32'b11111111111111111111111110100011;
reg [32-1:0] bias_reg_48 = 32'b00000000000000000000000001001101;
reg [32-1:0] bias_reg_49 = 32'b11111111111111111111111111010110;
reg [32-1:0] bias_reg_50 = 32'b00000000000000000000000011001111;
reg [32-1:0] bias_reg_51 = 32'b11111111111111111111111111110101;
reg [32-1:0] bias_reg_52 = 32'b00000000000000000000000010110100;
reg [32-1:0] bias_reg_53 = 32'b00000000000000000000000011011101;
reg [32-1:0] bias_reg_54 = 32'b00000000000000000000000100100111;
reg [32-1:0] bias_reg_55 = 32'b00000000000000000000000001001000;
reg [32-1:0] bias_reg_56 = 32'b11111111111111111111111011001001;
reg [32-1:0] bias_reg_57 = 32'b00000000000000000000000001010011;
reg [32-1:0] bias_reg_58 = 32'b11111111111111111111111101001111;
reg [32-1:0] bias_reg_59 = 32'b00000000000000000000000011001100;
reg [32-1:0] bias_reg_60 = 32'b11111111111111111111110100010110;
reg [32-1:0] bias_reg_61 = 32'b11111111111111111111111111110010;
reg [32-1:0] bias_reg_62 = 32'b11111111111111111111111110110111;
reg [32-1:0] bias_reg_63 = 32'b00000000000000000000000001110001;
assign bias_mem[0] = bias_reg_0;
assign bias_mem[1] = bias_reg_1;
assign bias_mem[2] = bias_reg_2;
assign bias_mem[3] = bias_reg_3;
assign bias_mem[4] = bias_reg_4;
assign bias_mem[5] = bias_reg_5;
assign bias_mem[6] = bias_reg_6;
assign bias_mem[7] = bias_reg_7;
assign bias_mem[8] = bias_reg_8;
assign bias_mem[9] = bias_reg_9;
assign bias_mem[10] = bias_reg_10;
assign bias_mem[11] = bias_reg_11;
assign bias_mem[12] = bias_reg_12;
assign bias_mem[13] = bias_reg_13;
assign bias_mem[14] = bias_reg_14;
assign bias_mem[15] = bias_reg_15;
assign bias_mem[16] = bias_reg_16;
assign bias_mem[17] = bias_reg_17;
assign bias_mem[18] = bias_reg_18;
assign bias_mem[19] = bias_reg_19;
assign bias_mem[20] = bias_reg_20;
assign bias_mem[21] = bias_reg_21;
assign bias_mem[22] = bias_reg_22;
assign bias_mem[23] = bias_reg_23;
assign bias_mem[24] = bias_reg_24;
assign bias_mem[25] = bias_reg_25;
assign bias_mem[26] = bias_reg_26;
assign bias_mem[27] = bias_reg_27;
assign bias_mem[28] = bias_reg_28;
assign bias_mem[29] = bias_reg_29;
assign bias_mem[30] = bias_reg_30;
assign bias_mem[31] = bias_reg_31;
assign bias_mem[32] = bias_reg_32;
assign bias_mem[33] = bias_reg_33;
assign bias_mem[34] = bias_reg_34;
assign bias_mem[35] = bias_reg_35;
assign bias_mem[36] = bias_reg_36;
assign bias_mem[37] = bias_reg_37;
assign bias_mem[38] = bias_reg_38;
assign bias_mem[39] = bias_reg_39;
assign bias_mem[40] = bias_reg_40;
assign bias_mem[41] = bias_reg_41;
assign bias_mem[42] = bias_reg_42;
assign bias_mem[43] = bias_reg_43;
assign bias_mem[44] = bias_reg_44;
assign bias_mem[45] = bias_reg_45;
assign bias_mem[46] = bias_reg_46;
assign bias_mem[47] = bias_reg_47;
assign bias_mem[48] = bias_reg_48;
assign bias_mem[49] = bias_reg_49;
assign bias_mem[50] = bias_reg_50;
assign bias_mem[51] = bias_reg_51;
assign bias_mem[52] = bias_reg_52;
assign bias_mem[53] = bias_reg_53;
assign bias_mem[54] = bias_reg_54;
assign bias_mem[55] = bias_reg_55;
assign bias_mem[56] = bias_reg_56;
assign bias_mem[57] = bias_reg_57;
assign bias_mem[58] = bias_reg_58;
assign bias_mem[59] = bias_reg_59;
assign bias_mem[60] = bias_reg_60;
assign bias_mem[61] = bias_reg_61;
assign bias_mem[62] = bias_reg_62;
assign bias_mem[63] = bias_reg_63;
endmodule
