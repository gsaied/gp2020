
module biasing_fire3_expand1 (
	output [32-1:0] bias_mem [0:64-1]
);

parameter [32-1:0] bias_parameter_0 = 32'b11111111111111111111111010111111;
parameter [32-1:0] bias_parameter_1 = 32'b00000000000000000000000100100010;
parameter [32-1:0] bias_parameter_2 = 32'b00000000000000000000001011001010;
parameter [32-1:0] bias_parameter_3 = 32'b00000000000000000000010010010001;
parameter [32-1:0] bias_parameter_4 = 32'b00000000000000000000000010011010;
parameter [32-1:0] bias_parameter_5 = 32'b11111111111111111111111101111110;
parameter [32-1:0] bias_parameter_6 = 32'b00000000000000000000001000011101;
parameter [32-1:0] bias_parameter_7 = 32'b00000000000000000000000100101000;
parameter [32-1:0] bias_parameter_8 = 32'b00000000000000000000000000111100;
parameter [32-1:0] bias_parameter_9 = 32'b00000000000000000000000101111101;
parameter [32-1:0] bias_parameter_10 = 32'b11111111111111111111110101111110;
parameter [32-1:0] bias_parameter_11 = 32'b00000000000000000000000000111010;
parameter [32-1:0] bias_parameter_12 = 32'b00000000000000000000001101011110;
parameter [32-1:0] bias_parameter_13 = 32'b00000000000000000000000110101110;
parameter [32-1:0] bias_parameter_14 = 32'b00000000000000000000000001000100;
parameter [32-1:0] bias_parameter_15 = 32'b00000000000000000000001000000011;
parameter [32-1:0] bias_parameter_16 = 32'b11111111111111111111111111110010;
parameter [32-1:0] bias_parameter_17 = 32'b00000000000000000000000000011111;
parameter [32-1:0] bias_parameter_18 = 32'b11111111111111111111111111101111;
parameter [32-1:0] bias_parameter_19 = 32'b00000000000000000000000000001000;
parameter [32-1:0] bias_parameter_20 = 32'b00000000000000000000000011110011;
parameter [32-1:0] bias_parameter_21 = 32'b00000000000000000000000101110000;
parameter [32-1:0] bias_parameter_22 = 32'b00000000000000000000000010000010;
parameter [32-1:0] bias_parameter_23 = 32'b00000000000000000000000010000000;
parameter [32-1:0] bias_parameter_24 = 32'b00000000000000000000010000111000;
parameter [32-1:0] bias_parameter_25 = 32'b00000000000000000000000011000000;
parameter [32-1:0] bias_parameter_26 = 32'b00000000000000000000000011011010;
parameter [32-1:0] bias_parameter_27 = 32'b00000000000000000000000010011100;
parameter [32-1:0] bias_parameter_28 = 32'b00000000000000000000000110000110;
parameter [32-1:0] bias_parameter_29 = 32'b00000000000000000000000010011001;
parameter [32-1:0] bias_parameter_30 = 32'b00000000000000000000001010000110;
parameter [32-1:0] bias_parameter_31 = 32'b00000000000000000000000001100010;
parameter [32-1:0] bias_parameter_32 = 32'b00000000000000000000000000000000;
parameter [32-1:0] bias_parameter_33 = 32'b00000000000000000000000011100000;
parameter [32-1:0] bias_parameter_34 = 32'b11111111111111111111111111011000;
parameter [32-1:0] bias_parameter_35 = 32'b11111111111111111111111110101100;
parameter [32-1:0] bias_parameter_36 = 32'b11111111111111111111111110101100;
parameter [32-1:0] bias_parameter_37 = 32'b00000000000000000000001110011101;
parameter [32-1:0] bias_parameter_38 = 32'b00000000000000000000000110111000;
parameter [32-1:0] bias_parameter_39 = 32'b00000000000000000000000011001101;
parameter [32-1:0] bias_parameter_40 = 32'b00000000000000000000000100001001;
parameter [32-1:0] bias_parameter_41 = 32'b00000000000000000000000000111010;
parameter [32-1:0] bias_parameter_42 = 32'b11111111111111111111111110001011;
parameter [32-1:0] bias_parameter_43 = 32'b11111111111111111111111110011000;
parameter [32-1:0] bias_parameter_44 = 32'b11111111111111111111111111010111;
parameter [32-1:0] bias_parameter_45 = 32'b00000000000000000000000011000100;
parameter [32-1:0] bias_parameter_46 = 32'b11111111111111111111111101011111;
parameter [32-1:0] bias_parameter_47 = 32'b00000000000000000000000011100010;
parameter [32-1:0] bias_parameter_48 = 32'b00000000000000000000000100110010;
parameter [32-1:0] bias_parameter_49 = 32'b00000000000000000000000100010011;
parameter [32-1:0] bias_parameter_50 = 32'b00000000000000000000000101111110;
parameter [32-1:0] bias_parameter_51 = 32'b00000000000000000000000010000101;
parameter [32-1:0] bias_parameter_52 = 32'b11111111111111111111111101111000;
parameter [32-1:0] bias_parameter_53 = 32'b00000000000000000000000110100000;
parameter [32-1:0] bias_parameter_54 = 32'b00000000000000000000000111000000;
parameter [32-1:0] bias_parameter_55 = 32'b11111111111111111111111111001001;
parameter [32-1:0] bias_parameter_56 = 32'b00000000000000000000001011000101;
parameter [32-1:0] bias_parameter_57 = 32'b11111111111111111111111101111100;
parameter [32-1:0] bias_parameter_58 = 32'b11111111111111111111111101101010;
parameter [32-1:0] bias_parameter_59 = 32'b11111111111111111111111111000110;
parameter [32-1:0] bias_parameter_60 = 32'b00000000000000000000001001100000;
parameter [32-1:0] bias_parameter_61 = 32'b00000000000000000000001001001100;
parameter [32-1:0] bias_parameter_62 = 32'b11111111111111111111111101001001;
parameter [32-1:0] bias_parameter_63 = 32'b00000000000000000000000000000000;
assign bias_mem[0] = bias_parameter_0;
assign bias_mem[1] = bias_parameter_1;
assign bias_mem[2] = bias_parameter_2;
assign bias_mem[3] = bias_parameter_3;
assign bias_mem[4] = bias_parameter_4;
assign bias_mem[5] = bias_parameter_5;
assign bias_mem[6] = bias_parameter_6;
assign bias_mem[7] = bias_parameter_7;
assign bias_mem[8] = bias_parameter_8;
assign bias_mem[9] = bias_parameter_9;
assign bias_mem[10] = bias_parameter_10;
assign bias_mem[11] = bias_parameter_11;
assign bias_mem[12] = bias_parameter_12;
assign bias_mem[13] = bias_parameter_13;
assign bias_mem[14] = bias_parameter_14;
assign bias_mem[15] = bias_parameter_15;
assign bias_mem[16] = bias_parameter_16;
assign bias_mem[17] = bias_parameter_17;
assign bias_mem[18] = bias_parameter_18;
assign bias_mem[19] = bias_parameter_19;
assign bias_mem[20] = bias_parameter_20;
assign bias_mem[21] = bias_parameter_21;
assign bias_mem[22] = bias_parameter_22;
assign bias_mem[23] = bias_parameter_23;
assign bias_mem[24] = bias_parameter_24;
assign bias_mem[25] = bias_parameter_25;
assign bias_mem[26] = bias_parameter_26;
assign bias_mem[27] = bias_parameter_27;
assign bias_mem[28] = bias_parameter_28;
assign bias_mem[29] = bias_parameter_29;
assign bias_mem[30] = bias_parameter_30;
assign bias_mem[31] = bias_parameter_31;
assign bias_mem[32] = bias_parameter_32;
assign bias_mem[33] = bias_parameter_33;
assign bias_mem[34] = bias_parameter_34;
assign bias_mem[35] = bias_parameter_35;
assign bias_mem[36] = bias_parameter_36;
assign bias_mem[37] = bias_parameter_37;
assign bias_mem[38] = bias_parameter_38;
assign bias_mem[39] = bias_parameter_39;
assign bias_mem[40] = bias_parameter_40;
assign bias_mem[41] = bias_parameter_41;
assign bias_mem[42] = bias_parameter_42;
assign bias_mem[43] = bias_parameter_43;
assign bias_mem[44] = bias_parameter_44;
assign bias_mem[45] = bias_parameter_45;
assign bias_mem[46] = bias_parameter_46;
assign bias_mem[47] = bias_parameter_47;
assign bias_mem[48] = bias_parameter_48;
assign bias_mem[49] = bias_parameter_49;
assign bias_mem[50] = bias_parameter_50;
assign bias_mem[51] = bias_parameter_51;
assign bias_mem[52] = bias_parameter_52;
assign bias_mem[53] = bias_parameter_53;
assign bias_mem[54] = bias_parameter_54;
assign bias_mem[55] = bias_parameter_55;
assign bias_mem[56] = bias_parameter_56;
assign bias_mem[57] = bias_parameter_57;
assign bias_mem[58] = bias_parameter_58;
assign bias_mem[59] = bias_parameter_59;
assign bias_mem[60] = bias_parameter_60;
assign bias_mem[61] = bias_parameter_61;
assign bias_mem[62] = bias_parameter_62;
assign bias_mem[63] = bias_parameter_63;
endmodule
