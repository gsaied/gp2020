
module biasing_fire9Squeeze (
	output [32-1:0] bias_mem [0:112-1]
);

reg [32-1:0] bias_reg_0 = 32'b00000000000000000000000110011110;
reg [32-1:0] bias_reg_1 = 32'b11111111111111111111110110100011;
reg [32-1:0] bias_reg_2 = 32'b00000000000000000000000101001011;
reg [32-1:0] bias_reg_3 = 32'b00000000000000000000000011101110;
reg [32-1:0] bias_reg_4 = 32'b11111111111111111111110001000001;
reg [32-1:0] bias_reg_5 = 32'b11111111111111111111111010111000;
reg [32-1:0] bias_reg_6 = 32'b00000000000000000000000111111110;
reg [32-1:0] bias_reg_7 = 32'b11111111111111111111101001111011;
reg [32-1:0] bias_reg_8 = 32'b11111111111111111111110111110110;
reg [32-1:0] bias_reg_9 = 32'b11111111111111111111111110010000;
reg [32-1:0] bias_reg_10 = 32'b00000000000000000000000011100001;
reg [32-1:0] bias_reg_11 = 32'b11111111111111111111111011011000;
reg [32-1:0] bias_reg_12 = 32'b11111111111111111111111101100010;
reg [32-1:0] bias_reg_13 = 32'b00000000000000000000000100101011;
reg [32-1:0] bias_reg_14 = 32'b11111111111111111111111011000110;
reg [32-1:0] bias_reg_15 = 32'b11111111111111111111111101110001;
reg [32-1:0] bias_reg_16 = 32'b00000000000000000000000011110000;
reg [32-1:0] bias_reg_17 = 32'b11111111111111111111111011000000;
reg [32-1:0] bias_reg_18 = 32'b00000000000000000000000100000011;
reg [32-1:0] bias_reg_19 = 32'b00000000000000000000000101000000;
reg [32-1:0] bias_reg_20 = 32'b00000000000000000000001000101101;
reg [32-1:0] bias_reg_21 = 32'b11111111111111111111001111010000;
reg [32-1:0] bias_reg_22 = 32'b11111111111111111111111001011011;
reg [32-1:0] bias_reg_23 = 32'b00000000000000000000000011110110;
reg [32-1:0] bias_reg_24 = 32'b00000000000000000000001010100101;
reg [32-1:0] bias_reg_25 = 32'b00000000000000000000001000010100;
reg [32-1:0] bias_reg_26 = 32'b11111111111111111111111100111001;
reg [32-1:0] bias_reg_27 = 32'b00000000000000000000000000100010;
reg [32-1:0] bias_reg_28 = 32'b00000000000000000000000000100100;
reg [32-1:0] bias_reg_29 = 32'b00000000000000000000000100110011;
reg [32-1:0] bias_reg_30 = 32'b11111111111111111111111010100001;
reg [32-1:0] bias_reg_31 = 32'b00000000000000000000000010000101;
reg [32-1:0] bias_reg_32 = 32'b11111111111111111111111101010001;
reg [32-1:0] bias_reg_33 = 32'b00000000000000000000000001100000;
reg [32-1:0] bias_reg_34 = 32'b11111111111111111111110101100001;
reg [32-1:0] bias_reg_35 = 32'b11111111111111111111110011101100;
reg [32-1:0] bias_reg_36 = 32'b11111111111111111111111000010010;
reg [32-1:0] bias_reg_37 = 32'b11111111111111111110100000000111;
reg [32-1:0] bias_reg_38 = 32'b11111111111111111111101101010011;
reg [32-1:0] bias_reg_39 = 32'b00000000000000000000000000000010;
reg [32-1:0] bias_reg_40 = 32'b11111111111111111111110011001100;
reg [32-1:0] bias_reg_41 = 32'b00000000000000000000000101000101;
reg [32-1:0] bias_reg_42 = 32'b00000000000000000000001010101010;
reg [32-1:0] bias_reg_43 = 32'b11111111111111111111110011111101;
reg [32-1:0] bias_reg_44 = 32'b00000000000000000000001101110100;
reg [32-1:0] bias_reg_45 = 32'b00000000000000000000000011011111;
reg [32-1:0] bias_reg_46 = 32'b00000000000000000000000001100000;
reg [32-1:0] bias_reg_47 = 32'b11111111111111111111111111010010;
reg [32-1:0] bias_reg_48 = 32'b11111111111111111111111010111010;
reg [32-1:0] bias_reg_49 = 32'b11111111111111111111111111100100;
reg [32-1:0] bias_reg_50 = 32'b11111111111111111111110101111100;
reg [32-1:0] bias_reg_51 = 32'b11111111111111111111110000010110;
reg [32-1:0] bias_reg_52 = 32'b11111111111111111111111100000011;
reg [32-1:0] bias_reg_53 = 32'b00000000000000000000000000001010;
reg [32-1:0] bias_reg_54 = 32'b11111111111111111111111110001001;
reg [32-1:0] bias_reg_55 = 32'b00000000000000000000000011000010;
reg [32-1:0] bias_reg_56 = 32'b00000000000000000000000001110110;
reg [32-1:0] bias_reg_57 = 32'b11111111111111111111110011111010;
reg [32-1:0] bias_reg_58 = 32'b00000000000000000001001000110011;
reg [32-1:0] bias_reg_59 = 32'b00000000000000000000000011101010;
reg [32-1:0] bias_reg_60 = 32'b00000000000000000000000001101111;
reg [32-1:0] bias_reg_61 = 32'b11111111111111111111111111000100;
reg [32-1:0] bias_reg_62 = 32'b00000000000000000000000011011101;
reg [32-1:0] bias_reg_63 = 32'b00000000000000000000000100100011;
reg [32-1:0] bias_reg_64 = 32'b00000000000000000000001000010100;
reg [32-1:0] bias_reg_65 = 32'b00000000000000000000000000001000;
reg [32-1:0] bias_reg_66 = 32'b00000000000000000000000011000100;
reg [32-1:0] bias_reg_67 = 32'b00000000000000000000000010000000;
reg [32-1:0] bias_reg_68 = 32'b00000000000000000000000110111111;
reg [32-1:0] bias_reg_69 = 32'b11111111111111111111101110000100;
reg [32-1:0] bias_reg_70 = 32'b00000000000000000000000001001110;
reg [32-1:0] bias_reg_71 = 32'b11111111111111111111100100101110;
reg [32-1:0] bias_reg_72 = 32'b00000000000000000000001001001101;
reg [32-1:0] bias_reg_73 = 32'b11111111111111111111111111001010;
reg [32-1:0] bias_reg_74 = 32'b11111111111111111111111110111011;
reg [32-1:0] bias_reg_75 = 32'b11111111111111111111101010111101;
reg [32-1:0] bias_reg_76 = 32'b11111111111111111111111100010010;
reg [32-1:0] bias_reg_77 = 32'b00000000000000000000001010001100;
reg [32-1:0] bias_reg_78 = 32'b11111111111111111111111001011001;
reg [32-1:0] bias_reg_79 = 32'b00000000000000000000000100000110;
reg [32-1:0] bias_reg_80 = 32'b00000000000000000000000101001000;
reg [32-1:0] bias_reg_81 = 32'b11111111111111111111111111110110;
reg [32-1:0] bias_reg_82 = 32'b11111111111111111111111011111001;
reg [32-1:0] bias_reg_83 = 32'b00000000000000000000000010101110;
reg [32-1:0] bias_reg_84 = 32'b11111111111111111111111111010001;
reg [32-1:0] bias_reg_85 = 32'b00000000000000000000000010000000;
reg [32-1:0] bias_reg_86 = 32'b11111111111111111111101000010010;
reg [32-1:0] bias_reg_87 = 32'b11111111111111111111111000000001;
reg [32-1:0] bias_reg_88 = 32'b00000000000000000000001000100011;
reg [32-1:0] bias_reg_89 = 32'b00000000000000000000000011000111;
reg [32-1:0] bias_reg_90 = 32'b00000000000000000000000000100101;
reg [32-1:0] bias_reg_91 = 32'b00000000000000000000000100000111;
reg [32-1:0] bias_reg_92 = 32'b00000000000000000000000111010100;
reg [32-1:0] bias_reg_93 = 32'b11111111111111111111110011111101;
reg [32-1:0] bias_reg_94 = 32'b11111111111111111111110111101100;
reg [32-1:0] bias_reg_95 = 32'b11111111111111111111111011010011;
reg [32-1:0] bias_reg_96 = 32'b11111111111111111111111101000101;
reg [32-1:0] bias_reg_97 = 32'b11111111111111111111111111011101;
reg [32-1:0] bias_reg_98 = 32'b11111111111111111111101011001001;
reg [32-1:0] bias_reg_99 = 32'b00000000000000000000000110111000;
reg [32-1:0] bias_reg_100 = 32'b11111111111111111111111101010111;
reg [32-1:0] bias_reg_101 = 32'b00000000000000000000000110011110;
reg [32-1:0] bias_reg_102 = 32'b00000000000000000000000100101100;
reg [32-1:0] bias_reg_103 = 32'b00000000000000000000001010000000;
reg [32-1:0] bias_reg_104 = 32'b00000000000000000000000011011100;
reg [32-1:0] bias_reg_105 = 32'b11111111111111111111101111101101;
reg [32-1:0] bias_reg_106 = 32'b00000000000000000000000111100010;
reg [32-1:0] bias_reg_107 = 32'b11111111111111111111100111111011;
reg [32-1:0] bias_reg_108 = 32'b11111111111111111111111100110101;
reg [32-1:0] bias_reg_109 = 32'b00000000000000000000000011110011;
reg [32-1:0] bias_reg_110 = 32'b11111111111111111111111110101001;
reg [32-1:0] bias_reg_111 = 32'b11111111111111111111111011000001;
assign bias_mem[0] = bias_reg_0;
assign bias_mem[1] = bias_reg_1;
assign bias_mem[2] = bias_reg_2;
assign bias_mem[3] = bias_reg_3;
assign bias_mem[4] = bias_reg_4;
assign bias_mem[5] = bias_reg_5;
assign bias_mem[6] = bias_reg_6;
assign bias_mem[7] = bias_reg_7;
assign bias_mem[8] = bias_reg_8;
assign bias_mem[9] = bias_reg_9;
assign bias_mem[10] = bias_reg_10;
assign bias_mem[11] = bias_reg_11;
assign bias_mem[12] = bias_reg_12;
assign bias_mem[13] = bias_reg_13;
assign bias_mem[14] = bias_reg_14;
assign bias_mem[15] = bias_reg_15;
assign bias_mem[16] = bias_reg_16;
assign bias_mem[17] = bias_reg_17;
assign bias_mem[18] = bias_reg_18;
assign bias_mem[19] = bias_reg_19;
assign bias_mem[20] = bias_reg_20;
assign bias_mem[21] = bias_reg_21;
assign bias_mem[22] = bias_reg_22;
assign bias_mem[23] = bias_reg_23;
assign bias_mem[24] = bias_reg_24;
assign bias_mem[25] = bias_reg_25;
assign bias_mem[26] = bias_reg_26;
assign bias_mem[27] = bias_reg_27;
assign bias_mem[28] = bias_reg_28;
assign bias_mem[29] = bias_reg_29;
assign bias_mem[30] = bias_reg_30;
assign bias_mem[31] = bias_reg_31;
assign bias_mem[32] = bias_reg_32;
assign bias_mem[33] = bias_reg_33;
assign bias_mem[34] = bias_reg_34;
assign bias_mem[35] = bias_reg_35;
assign bias_mem[36] = bias_reg_36;
assign bias_mem[37] = bias_reg_37;
assign bias_mem[38] = bias_reg_38;
assign bias_mem[39] = bias_reg_39;
assign bias_mem[40] = bias_reg_40;
assign bias_mem[41] = bias_reg_41;
assign bias_mem[42] = bias_reg_42;
assign bias_mem[43] = bias_reg_43;
assign bias_mem[44] = bias_reg_44;
assign bias_mem[45] = bias_reg_45;
assign bias_mem[46] = bias_reg_46;
assign bias_mem[47] = bias_reg_47;
assign bias_mem[48] = bias_reg_48;
assign bias_mem[49] = bias_reg_49;
assign bias_mem[50] = bias_reg_50;
assign bias_mem[51] = bias_reg_51;
assign bias_mem[52] = bias_reg_52;
assign bias_mem[53] = bias_reg_53;
assign bias_mem[54] = bias_reg_54;
assign bias_mem[55] = bias_reg_55;
assign bias_mem[56] = bias_reg_56;
assign bias_mem[57] = bias_reg_57;
assign bias_mem[58] = bias_reg_58;
assign bias_mem[59] = bias_reg_59;
assign bias_mem[60] = bias_reg_60;
assign bias_mem[61] = bias_reg_61;
assign bias_mem[62] = bias_reg_62;
assign bias_mem[63] = bias_reg_63;
assign bias_mem[64] = bias_reg_64;
assign bias_mem[65] = bias_reg_65;
assign bias_mem[66] = bias_reg_66;
assign bias_mem[67] = bias_reg_67;
assign bias_mem[68] = bias_reg_68;
assign bias_mem[69] = bias_reg_69;
assign bias_mem[70] = bias_reg_70;
assign bias_mem[71] = bias_reg_71;
assign bias_mem[72] = bias_reg_72;
assign bias_mem[73] = bias_reg_73;
assign bias_mem[74] = bias_reg_74;
assign bias_mem[75] = bias_reg_75;
assign bias_mem[76] = bias_reg_76;
assign bias_mem[77] = bias_reg_77;
assign bias_mem[78] = bias_reg_78;
assign bias_mem[79] = bias_reg_79;
assign bias_mem[80] = bias_reg_80;
assign bias_mem[81] = bias_reg_81;
assign bias_mem[82] = bias_reg_82;
assign bias_mem[83] = bias_reg_83;
assign bias_mem[84] = bias_reg_84;
assign bias_mem[85] = bias_reg_85;
assign bias_mem[86] = bias_reg_86;
assign bias_mem[87] = bias_reg_87;
assign bias_mem[88] = bias_reg_88;
assign bias_mem[89] = bias_reg_89;
assign bias_mem[90] = bias_reg_90;
assign bias_mem[91] = bias_reg_91;
assign bias_mem[92] = bias_reg_92;
assign bias_mem[93] = bias_reg_93;
assign bias_mem[94] = bias_reg_94;
assign bias_mem[95] = bias_reg_95;
assign bias_mem[96] = bias_reg_96;
assign bias_mem[97] = bias_reg_97;
assign bias_mem[98] = bias_reg_98;
assign bias_mem[99] = bias_reg_99;
assign bias_mem[100] = bias_reg_100;
assign bias_mem[101] = bias_reg_101;
assign bias_mem[102] = bias_reg_102;
assign bias_mem[103] = bias_reg_103;
assign bias_mem[104] = bias_reg_104;
assign bias_mem[105] = bias_reg_105;
assign bias_mem[106] = bias_reg_106;
assign bias_mem[107] = bias_reg_107;
assign bias_mem[108] = bias_reg_108;
assign bias_mem[109] = bias_reg_109;
assign bias_mem[110] = bias_reg_110;
assign bias_mem[111] = bias_reg_111;
endmodule
