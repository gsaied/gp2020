
module biasing_conv10_1 (
	output [32-1:0] bias_mem [0:512-1]
);

reg [32-1:0] bias_reg_0 = 32'b11111111111111111111111111010100;
reg [32-1:0] bias_reg_1 = 32'b00000000000000000000000011101111;
reg [32-1:0] bias_reg_2 = 32'b11111111111111111111111111100011;
reg [32-1:0] bias_reg_3 = 32'b11111111111111111111111010011101;
reg [32-1:0] bias_reg_4 = 32'b00000000000000000000000000110010;
reg [32-1:0] bias_reg_5 = 32'b11111111111111111111110111010011;
reg [32-1:0] bias_reg_6 = 32'b00000000000000000000000110111000;
reg [32-1:0] bias_reg_7 = 32'b11111111111111111111111101011011;
reg [32-1:0] bias_reg_8 = 32'b11111111111111111111111101001111;
reg [32-1:0] bias_reg_9 = 32'b11111111111111111111111101011000;
reg [32-1:0] bias_reg_10 = 32'b11111111111111111111111111000010;
reg [32-1:0] bias_reg_11 = 32'b11111111111111111111111110011101;
reg [32-1:0] bias_reg_12 = 32'b00000000000000000000000001111110;
reg [32-1:0] bias_reg_13 = 32'b00000000000000000000000000011101;
reg [32-1:0] bias_reg_14 = 32'b00000000000000000000000000001110;
reg [32-1:0] bias_reg_15 = 32'b11111111111111111111111110101100;
reg [32-1:0] bias_reg_16 = 32'b11111111111111111111111010110111;
reg [32-1:0] bias_reg_17 = 32'b11111111111111111111111100011011;
reg [32-1:0] bias_reg_18 = 32'b11111111111111111111111110001011;
reg [32-1:0] bias_reg_19 = 32'b11111111111111111111111110000111;
reg [32-1:0] bias_reg_20 = 32'b00000000000000000000000000100100;
reg [32-1:0] bias_reg_21 = 32'b00000000000000000000000001010010;
reg [32-1:0] bias_reg_22 = 32'b00000000000000000000000010010101;
reg [32-1:0] bias_reg_23 = 32'b00000000000000000000000000011111;
reg [32-1:0] bias_reg_24 = 32'b11111111111111111111111111010011;
reg [32-1:0] bias_reg_25 = 32'b00000000000000000000000010100001;
reg [32-1:0] bias_reg_26 = 32'b11111111111111111111111101001101;
reg [32-1:0] bias_reg_27 = 32'b00000000000000000000000001000011;
reg [32-1:0] bias_reg_28 = 32'b11111111111111111111111110110001;
reg [32-1:0] bias_reg_29 = 32'b00000000000000000000000000101110;
reg [32-1:0] bias_reg_30 = 32'b00000000000000000000000000011100;
reg [32-1:0] bias_reg_31 = 32'b00000000000000000000000001101110;
reg [32-1:0] bias_reg_32 = 32'b11111111111111111111111110101011;
reg [32-1:0] bias_reg_33 = 32'b11111111111111111111111010110010;
reg [32-1:0] bias_reg_34 = 32'b11111111111111111111111100011100;
reg [32-1:0] bias_reg_35 = 32'b11111111111111111111111011111100;
reg [32-1:0] bias_reg_36 = 32'b11111111111111111111111101111100;
reg [32-1:0] bias_reg_37 = 32'b00000000000000000000000011111110;
reg [32-1:0] bias_reg_38 = 32'b00000000000000000000000000101000;
reg [32-1:0] bias_reg_39 = 32'b11111111111111111111111011001100;
reg [32-1:0] bias_reg_40 = 32'b00000000000000000000000001111011;
reg [32-1:0] bias_reg_41 = 32'b11111111111111111111111111011100;
reg [32-1:0] bias_reg_42 = 32'b00000000000000000000000010110111;
reg [32-1:0] bias_reg_43 = 32'b11111111111111111111111100100110;
reg [32-1:0] bias_reg_44 = 32'b11111111111111111111111110101011;
reg [32-1:0] bias_reg_45 = 32'b00000000000000000000000101001000;
reg [32-1:0] bias_reg_46 = 32'b00000000000000000000000001011000;
reg [32-1:0] bias_reg_47 = 32'b11111111111111111111111010111011;
reg [32-1:0] bias_reg_48 = 32'b00000000000000000000000010111111;
reg [32-1:0] bias_reg_49 = 32'b00000000000000000000000010101101;
reg [32-1:0] bias_reg_50 = 32'b00000000000000000000000011100110;
reg [32-1:0] bias_reg_51 = 32'b11111111111111111111111110101000;
reg [32-1:0] bias_reg_52 = 32'b00000000000000000000000001011000;
reg [32-1:0] bias_reg_53 = 32'b00000000000000000000000000000111;
reg [32-1:0] bias_reg_54 = 32'b11111111111111111111111110001001;
reg [32-1:0] bias_reg_55 = 32'b11111111111111111111111111010000;
reg [32-1:0] bias_reg_56 = 32'b00000000000000000000000010101001;
reg [32-1:0] bias_reg_57 = 32'b00000000000000000000000010110101;
reg [32-1:0] bias_reg_58 = 32'b00000000000000000000001101110000;
reg [32-1:0] bias_reg_59 = 32'b00000000000000000000000000001011;
reg [32-1:0] bias_reg_60 = 32'b11111111111111111111111100010101;
reg [32-1:0] bias_reg_61 = 32'b00000000000000000000000110001001;
reg [32-1:0] bias_reg_62 = 32'b11111111111111111111111011111111;
reg [32-1:0] bias_reg_63 = 32'b00000000000000000000000001000010;
reg [32-1:0] bias_reg_64 = 32'b00000000000000000000000100100110;
reg [32-1:0] bias_reg_65 = 32'b00000000000000000000000000100111;
reg [32-1:0] bias_reg_66 = 32'b11111111111111111111111100101001;
reg [32-1:0] bias_reg_67 = 32'b11111111111111111111111101101101;
reg [32-1:0] bias_reg_68 = 32'b11111111111111111111111011101101;
reg [32-1:0] bias_reg_69 = 32'b00000000000000000000000100000111;
reg [32-1:0] bias_reg_70 = 32'b00000000000000000000000000111111;
reg [32-1:0] bias_reg_71 = 32'b11111111111111111111111101010000;
reg [32-1:0] bias_reg_72 = 32'b11111111111111111111111110001100;
reg [32-1:0] bias_reg_73 = 32'b11111111111111111111111011011101;
reg [32-1:0] bias_reg_74 = 32'b00000000000000000000000000000001;
reg [32-1:0] bias_reg_75 = 32'b00000000000000000000000001110010;
reg [32-1:0] bias_reg_76 = 32'b00000000000000000000000000010101;
reg [32-1:0] bias_reg_77 = 32'b00000000000000000000000101010101;
reg [32-1:0] bias_reg_78 = 32'b11111111111111111111111011000111;
reg [32-1:0] bias_reg_79 = 32'b00000000000000000000000011011001;
reg [32-1:0] bias_reg_80 = 32'b11111111111111111111111001111111;
reg [32-1:0] bias_reg_81 = 32'b11111111111111111111111101010101;
reg [32-1:0] bias_reg_82 = 32'b11111111111111111111111110101001;
reg [32-1:0] bias_reg_83 = 32'b11111111111111111111111101010000;
reg [32-1:0] bias_reg_84 = 32'b11111111111111111111111010001100;
reg [32-1:0] bias_reg_85 = 32'b11111111111111111111111111000110;
reg [32-1:0] bias_reg_86 = 32'b11111111111111111111111101100000;
reg [32-1:0] bias_reg_87 = 32'b11111111111111111111111110010110;
reg [32-1:0] bias_reg_88 = 32'b11111111111111111111111110011111;
reg [32-1:0] bias_reg_89 = 32'b00000000000000000000000010010001;
reg [32-1:0] bias_reg_90 = 32'b11111111111111111111111101101111;
reg [32-1:0] bias_reg_91 = 32'b00000000000000000000000000100101;
reg [32-1:0] bias_reg_92 = 32'b00000000000000000000000000111010;
reg [32-1:0] bias_reg_93 = 32'b11111111111111111111111101110011;
reg [32-1:0] bias_reg_94 = 32'b00000000000000000000000001101010;
reg [32-1:0] bias_reg_95 = 32'b00000000000000000000000000000100;
reg [32-1:0] bias_reg_96 = 32'b00000000000000000000000010010011;
reg [32-1:0] bias_reg_97 = 32'b11111111111111111111111111100111;
reg [32-1:0] bias_reg_98 = 32'b11111111111111111111111100011000;
reg [32-1:0] bias_reg_99 = 32'b11111111111111111111111100011010;
reg [32-1:0] bias_reg_100 = 32'b11111111111111111111111011111011;
reg [32-1:0] bias_reg_101 = 32'b11111111111111111111111001111000;
reg [32-1:0] bias_reg_102 = 32'b00000000000000000000000011010101;
reg [32-1:0] bias_reg_103 = 32'b00000000000000000000000110100011;
reg [32-1:0] bias_reg_104 = 32'b00000000000000000000000010010100;
reg [32-1:0] bias_reg_105 = 32'b11111111111111111111111100000101;
reg [32-1:0] bias_reg_106 = 32'b00000000000000000000000011110111;
reg [32-1:0] bias_reg_107 = 32'b11111111111111111111111101101101;
reg [32-1:0] bias_reg_108 = 32'b00000000000000000000000010111111;
reg [32-1:0] bias_reg_109 = 32'b00000000000000000000000000001111;
reg [32-1:0] bias_reg_110 = 32'b11111111111111111111111110000110;
reg [32-1:0] bias_reg_111 = 32'b00000000000000000000000111010110;
reg [32-1:0] bias_reg_112 = 32'b00000000000000000000000001111101;
reg [32-1:0] bias_reg_113 = 32'b00000000000000000000000001000001;
reg [32-1:0] bias_reg_114 = 32'b00000000000000000000000000100000;
reg [32-1:0] bias_reg_115 = 32'b00000000000000000000000001011101;
reg [32-1:0] bias_reg_116 = 32'b00000000000000000000000100100000;
reg [32-1:0] bias_reg_117 = 32'b11111111111111111111111101100111;
reg [32-1:0] bias_reg_118 = 32'b00000000000000000000000001011000;
reg [32-1:0] bias_reg_119 = 32'b00000000000000000000000001010101;
reg [32-1:0] bias_reg_120 = 32'b00000000000000000000000010110110;
reg [32-1:0] bias_reg_121 = 32'b11111111111111111111111101000111;
reg [32-1:0] bias_reg_122 = 32'b00000000000000000000000010001010;
reg [32-1:0] bias_reg_123 = 32'b11111111111111111111111110000100;
reg [32-1:0] bias_reg_124 = 32'b00000000000000000000000000001011;
reg [32-1:0] bias_reg_125 = 32'b00000000000000000000000000111000;
reg [32-1:0] bias_reg_126 = 32'b11111111111111111111110111101110;
reg [32-1:0] bias_reg_127 = 32'b11111111111111111111111100101001;
reg [32-1:0] bias_reg_128 = 32'b11111111111111111111111100110110;
reg [32-1:0] bias_reg_129 = 32'b00000000000000000000000100001111;
reg [32-1:0] bias_reg_130 = 32'b11111111111111111111111111100011;
reg [32-1:0] bias_reg_131 = 32'b11111111111111111111111010111110;
reg [32-1:0] bias_reg_132 = 32'b11111111111111111111111101111000;
reg [32-1:0] bias_reg_133 = 32'b00000000000000000000000010110101;
reg [32-1:0] bias_reg_134 = 32'b11111111111111111111111001011001;
reg [32-1:0] bias_reg_135 = 32'b11111111111111111111111110010111;
reg [32-1:0] bias_reg_136 = 32'b11111111111111111111111100010001;
reg [32-1:0] bias_reg_137 = 32'b11111111111111111111111111101100;
reg [32-1:0] bias_reg_138 = 32'b00000000000000000000000000001111;
reg [32-1:0] bias_reg_139 = 32'b00000000000000000000000000000111;
reg [32-1:0] bias_reg_140 = 32'b11111111111111111111111101010100;
reg [32-1:0] bias_reg_141 = 32'b11111111111111111111111111000000;
reg [32-1:0] bias_reg_142 = 32'b00000000000000000000000011100011;
reg [32-1:0] bias_reg_143 = 32'b11111111111111111111111110100011;
reg [32-1:0] bias_reg_144 = 32'b11111111111111111111111100010000;
reg [32-1:0] bias_reg_145 = 32'b11111111111111111111111110010100;
reg [32-1:0] bias_reg_146 = 32'b11111111111111111111111101011001;
reg [32-1:0] bias_reg_147 = 32'b11111111111111111111111101011110;
reg [32-1:0] bias_reg_148 = 32'b11111111111111111111111011000000;
reg [32-1:0] bias_reg_149 = 32'b00000000000000000000000001001000;
reg [32-1:0] bias_reg_150 = 32'b11111111111111111111111111110000;
reg [32-1:0] bias_reg_151 = 32'b00000000000000000000000000001101;
reg [32-1:0] bias_reg_152 = 32'b11111111111111111111111011000111;
reg [32-1:0] bias_reg_153 = 32'b00000000000000000000000001001110;
reg [32-1:0] bias_reg_154 = 32'b11111111111111111111111111000000;
reg [32-1:0] bias_reg_155 = 32'b11111111111111111111111110100100;
reg [32-1:0] bias_reg_156 = 32'b00000000000000000000000000101111;
reg [32-1:0] bias_reg_157 = 32'b11111111111111111111111100100111;
reg [32-1:0] bias_reg_158 = 32'b11111111111111111111111000010000;
reg [32-1:0] bias_reg_159 = 32'b11111111111111111111111111011110;
reg [32-1:0] bias_reg_160 = 32'b11111111111111111111111101111001;
reg [32-1:0] bias_reg_161 = 32'b00000000000000000000000010001011;
reg [32-1:0] bias_reg_162 = 32'b00000000000000000000000011011100;
reg [32-1:0] bias_reg_163 = 32'b11111111111111111111111111001101;
reg [32-1:0] bias_reg_164 = 32'b11111111111111111111111101111110;
reg [32-1:0] bias_reg_165 = 32'b11111111111111111111111110011001;
reg [32-1:0] bias_reg_166 = 32'b11111111111111111111111110110100;
reg [32-1:0] bias_reg_167 = 32'b11111111111111111111111101101100;
reg [32-1:0] bias_reg_168 = 32'b11111111111111111111111011001011;
reg [32-1:0] bias_reg_169 = 32'b00000000000000000000000001010100;
reg [32-1:0] bias_reg_170 = 32'b11111111111111111111111100110100;
reg [32-1:0] bias_reg_171 = 32'b00000000000000000000000000110111;
reg [32-1:0] bias_reg_172 = 32'b00000000000000000000000000111010;
reg [32-1:0] bias_reg_173 = 32'b00000000000000000000000001001101;
reg [32-1:0] bias_reg_174 = 32'b00000000000000000000000000011000;
reg [32-1:0] bias_reg_175 = 32'b11111111111111111111111101001111;
reg [32-1:0] bias_reg_176 = 32'b11111111111111111111110110111101;
reg [32-1:0] bias_reg_177 = 32'b11111111111111111111111111001110;
reg [32-1:0] bias_reg_178 = 32'b11111111111111111111111110100110;
reg [32-1:0] bias_reg_179 = 32'b11111111111111111111111110110000;
reg [32-1:0] bias_reg_180 = 32'b11111111111111111111111011000011;
reg [32-1:0] bias_reg_181 = 32'b11111111111111111111111110011100;
reg [32-1:0] bias_reg_182 = 32'b11111111111111111111111110000000;
reg [32-1:0] bias_reg_183 = 32'b00000000000000000000000010110100;
reg [32-1:0] bias_reg_184 = 32'b00000000000000000000000001000110;
reg [32-1:0] bias_reg_185 = 32'b00000000000000000000000001010001;
reg [32-1:0] bias_reg_186 = 32'b11111111111111111111111110001101;
reg [32-1:0] bias_reg_187 = 32'b00000000000000000000000001001011;
reg [32-1:0] bias_reg_188 = 32'b11111111111111111111111111110010;
reg [32-1:0] bias_reg_189 = 32'b11111111111111111111110111100101;
reg [32-1:0] bias_reg_190 = 32'b11111111111111111111111110110111;
reg [32-1:0] bias_reg_191 = 32'b11111111111111111111111100100101;
reg [32-1:0] bias_reg_192 = 32'b00000000000000000000000000000100;
reg [32-1:0] bias_reg_193 = 32'b11111111111111111111111000011010;
reg [32-1:0] bias_reg_194 = 32'b11111111111111111111111011001110;
reg [32-1:0] bias_reg_195 = 32'b00000000000000000000000001011010;
reg [32-1:0] bias_reg_196 = 32'b11111111111111111111111101111111;
reg [32-1:0] bias_reg_197 = 32'b11111111111111111111111010001001;
reg [32-1:0] bias_reg_198 = 32'b11111111111111111111111001100111;
reg [32-1:0] bias_reg_199 = 32'b00000000000000000000000001110100;
reg [32-1:0] bias_reg_200 = 32'b11111111111111111111111011101011;
reg [32-1:0] bias_reg_201 = 32'b11111111111111111111111101001010;
reg [32-1:0] bias_reg_202 = 32'b00000000000000000000000111111010;
reg [32-1:0] bias_reg_203 = 32'b00000000000000000000000010011010;
reg [32-1:0] bias_reg_204 = 32'b11111111111111111111111001001100;
reg [32-1:0] bias_reg_205 = 32'b11111111111111111111111100111000;
reg [32-1:0] bias_reg_206 = 32'b11111111111111111111111100001000;
reg [32-1:0] bias_reg_207 = 32'b11111111111111111111111101001000;
reg [32-1:0] bias_reg_208 = 32'b11111111111111111111111010111010;
reg [32-1:0] bias_reg_209 = 32'b00000000000000000000000101101111;
reg [32-1:0] bias_reg_210 = 32'b11111111111111111111111111100010;
reg [32-1:0] bias_reg_211 = 32'b00000000000000000000000111101000;
reg [32-1:0] bias_reg_212 = 32'b11111111111111111111111100001101;
reg [32-1:0] bias_reg_213 = 32'b00000000000000000000000100010110;
reg [32-1:0] bias_reg_214 = 32'b11111111111111111111111111001010;
reg [32-1:0] bias_reg_215 = 32'b00000000000000000000000010100001;
reg [32-1:0] bias_reg_216 = 32'b11111111111111111111111111001110;
reg [32-1:0] bias_reg_217 = 32'b00000000000000000000001000001011;
reg [32-1:0] bias_reg_218 = 32'b00000000000000000000000000011010;
reg [32-1:0] bias_reg_219 = 32'b11111111111111111111111111111111;
reg [32-1:0] bias_reg_220 = 32'b11111111111111111111111101001100;
reg [32-1:0] bias_reg_221 = 32'b00000000000000000000000001010111;
reg [32-1:0] bias_reg_222 = 32'b11111111111111111111111101111100;
reg [32-1:0] bias_reg_223 = 32'b00000000000000000000000101110100;
reg [32-1:0] bias_reg_224 = 32'b11111111111111111111111100100000;
reg [32-1:0] bias_reg_225 = 32'b00000000000000000000000001001001;
reg [32-1:0] bias_reg_226 = 32'b11111111111111111111111111101011;
reg [32-1:0] bias_reg_227 = 32'b11111111111111111111111100000011;
reg [32-1:0] bias_reg_228 = 32'b11111111111111111111111110011100;
reg [32-1:0] bias_reg_229 = 32'b00000000000000000000000011110010;
reg [32-1:0] bias_reg_230 = 32'b11111111111111111111111111111100;
reg [32-1:0] bias_reg_231 = 32'b11111111111111111111111010111000;
reg [32-1:0] bias_reg_232 = 32'b00000000000000000000000001111101;
reg [32-1:0] bias_reg_233 = 32'b11111111111111111111111011001011;
reg [32-1:0] bias_reg_234 = 32'b00000000000000000000000001011100;
reg [32-1:0] bias_reg_235 = 32'b11111111111111111111111101101100;
reg [32-1:0] bias_reg_236 = 32'b11111111111111111111111101011001;
reg [32-1:0] bias_reg_237 = 32'b00000000000000000000001000011011;
reg [32-1:0] bias_reg_238 = 32'b11111111111111111111111111011011;
reg [32-1:0] bias_reg_239 = 32'b00000000000000000000000010101000;
reg [32-1:0] bias_reg_240 = 32'b11111111111111111111111001110101;
reg [32-1:0] bias_reg_241 = 32'b00000000000000000000000001110010;
reg [32-1:0] bias_reg_242 = 32'b11111111111111111111111101111101;
reg [32-1:0] bias_reg_243 = 32'b11111111111111111111111101111011;
reg [32-1:0] bias_reg_244 = 32'b11111111111111111111111001101010;
reg [32-1:0] bias_reg_245 = 32'b11111111111111111111111110111001;
reg [32-1:0] bias_reg_246 = 32'b11111111111111111111111010100110;
reg [32-1:0] bias_reg_247 = 32'b11111111111111111111111111001100;
reg [32-1:0] bias_reg_248 = 32'b11111111111111111111111000101110;
reg [32-1:0] bias_reg_249 = 32'b11111111111111111111111101000100;
reg [32-1:0] bias_reg_250 = 32'b11111111111111111111111100000100;
reg [32-1:0] bias_reg_251 = 32'b00000000000000000000000000010110;
reg [32-1:0] bias_reg_252 = 32'b11111111111111111111111110101000;
reg [32-1:0] bias_reg_253 = 32'b11111111111111111111111100110001;
reg [32-1:0] bias_reg_254 = 32'b11111111111111111111111111100110;
reg [32-1:0] bias_reg_255 = 32'b11111111111111111111111101001011;
reg [32-1:0] bias_reg_256 = 32'b11111111111111111111111100000111;
reg [32-1:0] bias_reg_257 = 32'b11111111111111111111111111010101;
reg [32-1:0] bias_reg_258 = 32'b00000000000000000000000001111001;
reg [32-1:0] bias_reg_259 = 32'b11111111111111111111111101101011;
reg [32-1:0] bias_reg_260 = 32'b11111111111111111111111110000101;
reg [32-1:0] bias_reg_261 = 32'b00000000000000000000000001110111;
reg [32-1:0] bias_reg_262 = 32'b11111111111111111111111101000111;
reg [32-1:0] bias_reg_263 = 32'b00000000000000000000000100010101;
reg [32-1:0] bias_reg_264 = 32'b11111111111111111111111101111101;
reg [32-1:0] bias_reg_265 = 32'b11111111111111111111111000100110;
reg [32-1:0] bias_reg_266 = 32'b11111111111111111111111111100111;
reg [32-1:0] bias_reg_267 = 32'b11111111111111111111111010000111;
reg [32-1:0] bias_reg_268 = 32'b11111111111111111111111101100101;
reg [32-1:0] bias_reg_269 = 32'b11111111111111111111111101100000;
reg [32-1:0] bias_reg_270 = 32'b00000000000000000000000000110101;
reg [32-1:0] bias_reg_271 = 32'b11111111111111111111111100000000;
reg [32-1:0] bias_reg_272 = 32'b00000000000000000000000001010100;
reg [32-1:0] bias_reg_273 = 32'b00000000000000000000000101110111;
reg [32-1:0] bias_reg_274 = 32'b00000000000000000000000000111110;
reg [32-1:0] bias_reg_275 = 32'b00000000000000000000000001001101;
reg [32-1:0] bias_reg_276 = 32'b00000000000000000000000001001000;
reg [32-1:0] bias_reg_277 = 32'b00000000000000000000000001001000;
reg [32-1:0] bias_reg_278 = 32'b11111111111111111111111111111110;
reg [32-1:0] bias_reg_279 = 32'b11111111111111111111111100100000;
reg [32-1:0] bias_reg_280 = 32'b11111111111111111111111010111010;
reg [32-1:0] bias_reg_281 = 32'b00000000000000000000000100110010;
reg [32-1:0] bias_reg_282 = 32'b11111111111111111111111010100100;
reg [32-1:0] bias_reg_283 = 32'b00000000000000000000000000101110;
reg [32-1:0] bias_reg_284 = 32'b00000000000000000000000100010001;
reg [32-1:0] bias_reg_285 = 32'b00000000000000000000000000011010;
reg [32-1:0] bias_reg_286 = 32'b00000000000000000000000010011011;
reg [32-1:0] bias_reg_287 = 32'b11111111111111111111111111101100;
reg [32-1:0] bias_reg_288 = 32'b11111111111111111111111010001001;
reg [32-1:0] bias_reg_289 = 32'b00000000000000000000000010001010;
reg [32-1:0] bias_reg_290 = 32'b00000000000000000000000001110000;
reg [32-1:0] bias_reg_291 = 32'b00000000000000000000000001011011;
reg [32-1:0] bias_reg_292 = 32'b00000000000000000000000000101011;
reg [32-1:0] bias_reg_293 = 32'b11111111111111111111111101011100;
reg [32-1:0] bias_reg_294 = 32'b00000000000000000000000000011110;
reg [32-1:0] bias_reg_295 = 32'b00000000000000000000000100111011;
reg [32-1:0] bias_reg_296 = 32'b11111111111111111111111100100100;
reg [32-1:0] bias_reg_297 = 32'b00000000000000000000000000011011;
reg [32-1:0] bias_reg_298 = 32'b11111111111111111111111111010000;
reg [32-1:0] bias_reg_299 = 32'b00000000000000000000000011011001;
reg [32-1:0] bias_reg_300 = 32'b11111111111111111111111110011011;
reg [32-1:0] bias_reg_301 = 32'b00000000000000000000000000111000;
reg [32-1:0] bias_reg_302 = 32'b11111111111111111111111001100000;
reg [32-1:0] bias_reg_303 = 32'b11111111111111111111111011010011;
reg [32-1:0] bias_reg_304 = 32'b11111111111111111111111101101011;
reg [32-1:0] bias_reg_305 = 32'b00000000000000000000000100111001;
reg [32-1:0] bias_reg_306 = 32'b00000000000000000000000001100111;
reg [32-1:0] bias_reg_307 = 32'b00000000000000000000000000101100;
reg [32-1:0] bias_reg_308 = 32'b11111111111111111111111001110100;
reg [32-1:0] bias_reg_309 = 32'b00000000000000000000000100000100;
reg [32-1:0] bias_reg_310 = 32'b00000000000000000000000001110001;
reg [32-1:0] bias_reg_311 = 32'b00000000000000000000000001000111;
reg [32-1:0] bias_reg_312 = 32'b00000000000000000000000010010101;
reg [32-1:0] bias_reg_313 = 32'b00000000000000000000010011110010;
reg [32-1:0] bias_reg_314 = 32'b00000000000000000000000110001110;
reg [32-1:0] bias_reg_315 = 32'b00000000000000000000000111011011;
reg [32-1:0] bias_reg_316 = 32'b11111111111111111111111111011010;
reg [32-1:0] bias_reg_317 = 32'b00000000000000000000000111001110;
reg [32-1:0] bias_reg_318 = 32'b00000000000000000000000000110010;
reg [32-1:0] bias_reg_319 = 32'b11111111111111111111111011100001;
reg [32-1:0] bias_reg_320 = 32'b11111111111111111111111111100011;
reg [32-1:0] bias_reg_321 = 32'b11111111111111111111111101100101;
reg [32-1:0] bias_reg_322 = 32'b11111111111111111111111100101101;
reg [32-1:0] bias_reg_323 = 32'b11111111111111111111111110101101;
reg [32-1:0] bias_reg_324 = 32'b11111111111111111111111111111000;
reg [32-1:0] bias_reg_325 = 32'b00000000000000000000000000011010;
reg [32-1:0] bias_reg_326 = 32'b11111111111111111111111100110000;
reg [32-1:0] bias_reg_327 = 32'b00000000000000000000000000001001;
reg [32-1:0] bias_reg_328 = 32'b11111111111111111111111111110110;
reg [32-1:0] bias_reg_329 = 32'b00000000000000000000000110001011;
reg [32-1:0] bias_reg_330 = 32'b00000000000000000000000001000100;
reg [32-1:0] bias_reg_331 = 32'b11111111111111111111111100010001;
reg [32-1:0] bias_reg_332 = 32'b00000000000000000000000001001100;
reg [32-1:0] bias_reg_333 = 32'b00000000000000000000000001101010;
reg [32-1:0] bias_reg_334 = 32'b11111111111111111111111100001101;
reg [32-1:0] bias_reg_335 = 32'b00000000000000000000000010001000;
reg [32-1:0] bias_reg_336 = 32'b00000000000000000000000111010001;
reg [32-1:0] bias_reg_337 = 32'b11111111111111111111111010101010;
reg [32-1:0] bias_reg_338 = 32'b11111111111111111111111111110110;
reg [32-1:0] bias_reg_339 = 32'b00000000000000000000001000010000;
reg [32-1:0] bias_reg_340 = 32'b11111111111111111111111110011000;
reg [32-1:0] bias_reg_341 = 32'b11111111111111111111111100001011;
reg [32-1:0] bias_reg_342 = 32'b11111111111111111111111011010100;
reg [32-1:0] bias_reg_343 = 32'b00000000000000000000000001010101;
reg [32-1:0] bias_reg_344 = 32'b00000000000000000000000010110101;
reg [32-1:0] bias_reg_345 = 32'b11111111111111111111111101111000;
reg [32-1:0] bias_reg_346 = 32'b00000000000000000000000011000110;
reg [32-1:0] bias_reg_347 = 32'b00000000000000000000000001101110;
reg [32-1:0] bias_reg_348 = 32'b11111111111111111111111110010100;
reg [32-1:0] bias_reg_349 = 32'b00000000000000000000000001001110;
reg [32-1:0] bias_reg_350 = 32'b11111111111111111111111111001011;
reg [32-1:0] bias_reg_351 = 32'b00000000000000000000000011111010;
reg [32-1:0] bias_reg_352 = 32'b11111111111111111111111110110001;
reg [32-1:0] bias_reg_353 = 32'b11111111111111111111111101010101;
reg [32-1:0] bias_reg_354 = 32'b00000000000000000000000001001111;
reg [32-1:0] bias_reg_355 = 32'b11111111111111111111111101100111;
reg [32-1:0] bias_reg_356 = 32'b11111111111111111111111010000010;
reg [32-1:0] bias_reg_357 = 32'b11111111111111111111111110001011;
reg [32-1:0] bias_reg_358 = 32'b00000000000000000000000000010101;
reg [32-1:0] bias_reg_359 = 32'b00000000000000000000000001101111;
reg [32-1:0] bias_reg_360 = 32'b11111111111111111111111110001011;
reg [32-1:0] bias_reg_361 = 32'b00000000000000000000000000111000;
reg [32-1:0] bias_reg_362 = 32'b11111111111111111111111111100001;
reg [32-1:0] bias_reg_363 = 32'b00000000000000000000000000010001;
reg [32-1:0] bias_reg_364 = 32'b00000000000000000000001000100000;
reg [32-1:0] bias_reg_365 = 32'b00000000000000000000000001101110;
reg [32-1:0] bias_reg_366 = 32'b11111111111111111111111110000001;
reg [32-1:0] bias_reg_367 = 32'b00000000000000000000000001001001;
reg [32-1:0] bias_reg_368 = 32'b11111111111111111111111100101001;
reg [32-1:0] bias_reg_369 = 32'b11111111111111111111111111100011;
reg [32-1:0] bias_reg_370 = 32'b11111111111111111111111100001110;
reg [32-1:0] bias_reg_371 = 32'b11111111111111111111111010001100;
reg [32-1:0] bias_reg_372 = 32'b11111111111111111111111111100101;
reg [32-1:0] bias_reg_373 = 32'b00000000000000000000000000001110;
reg [32-1:0] bias_reg_374 = 32'b11111111111111111111111101100101;
reg [32-1:0] bias_reg_375 = 32'b11111111111111111111111100010111;
reg [32-1:0] bias_reg_376 = 32'b00000000000000000000000010011011;
reg [32-1:0] bias_reg_377 = 32'b00000000000000000000000010100110;
reg [32-1:0] bias_reg_378 = 32'b00000000000000000000000011111010;
reg [32-1:0] bias_reg_379 = 32'b00000000000000000000000100101011;
reg [32-1:0] bias_reg_380 = 32'b11111111111111111111110010101100;
reg [32-1:0] bias_reg_381 = 32'b11111111111111111111111111110010;
reg [32-1:0] bias_reg_382 = 32'b00000000000000000000000100000111;
reg [32-1:0] bias_reg_383 = 32'b11111111111111111111111111010101;
reg [32-1:0] bias_reg_384 = 32'b11111111111111111111111100011100;
reg [32-1:0] bias_reg_385 = 32'b11111111111111111111111111000101;
reg [32-1:0] bias_reg_386 = 32'b00000000000000000000000001011110;
reg [32-1:0] bias_reg_387 = 32'b00000000000000000000000010010010;
reg [32-1:0] bias_reg_388 = 32'b00000000000000000000000001001110;
reg [32-1:0] bias_reg_389 = 32'b11111111111111111111111011011001;
reg [32-1:0] bias_reg_390 = 32'b11111111111111111111111001010111;
reg [32-1:0] bias_reg_391 = 32'b00000000000000000000000001001100;
reg [32-1:0] bias_reg_392 = 32'b11111111111111111111111011100011;
reg [32-1:0] bias_reg_393 = 32'b00000000000000000000000000010000;
reg [32-1:0] bias_reg_394 = 32'b11111111111111111111111010001101;
reg [32-1:0] bias_reg_395 = 32'b11111111111111111111111101000100;
reg [32-1:0] bias_reg_396 = 32'b11111111111111111111111111010111;
reg [32-1:0] bias_reg_397 = 32'b11111111111111111111111100101100;
reg [32-1:0] bias_reg_398 = 32'b11111111111111111111111110110001;
reg [32-1:0] bias_reg_399 = 32'b00000000000000000000000011001000;
reg [32-1:0] bias_reg_400 = 32'b11111111111111111111111111010101;
reg [32-1:0] bias_reg_401 = 32'b11111111111111111111111110001110;
reg [32-1:0] bias_reg_402 = 32'b11111111111111111111111110011010;
reg [32-1:0] bias_reg_403 = 32'b11111111111111111111111011000111;
reg [32-1:0] bias_reg_404 = 32'b11111111111111111111111110100110;
reg [32-1:0] bias_reg_405 = 32'b00000000000000000000000100011100;
reg [32-1:0] bias_reg_406 = 32'b00000000000000000000000010100101;
reg [32-1:0] bias_reg_407 = 32'b00000000000000000000000000011000;
reg [32-1:0] bias_reg_408 = 32'b11111111111111111111110100010001;
reg [32-1:0] bias_reg_409 = 32'b11111111111111111111110111101011;
reg [32-1:0] bias_reg_410 = 32'b00000000000000000000000111111011;
reg [32-1:0] bias_reg_411 = 32'b00000000000000000000000100101010;
reg [32-1:0] bias_reg_412 = 32'b11111111111111111111110100111101;
reg [32-1:0] bias_reg_413 = 32'b11111111111111111111111100010110;
reg [32-1:0] bias_reg_414 = 32'b00000000000000000000000011001011;
reg [32-1:0] bias_reg_415 = 32'b00000000000000000000000001010000;
reg [32-1:0] bias_reg_416 = 32'b00000000000000000000000111000101;
reg [32-1:0] bias_reg_417 = 32'b00000000000000000000000000000100;
reg [32-1:0] bias_reg_418 = 32'b11111111111111111111111110001110;
reg [32-1:0] bias_reg_419 = 32'b00000000000000000000000101010010;
reg [32-1:0] bias_reg_420 = 32'b11111111111111111111111011111110;
reg [32-1:0] bias_reg_421 = 32'b00000000000000000000000111111110;
reg [32-1:0] bias_reg_422 = 32'b11111111111111111111111011100110;
reg [32-1:0] bias_reg_423 = 32'b00000000000000000000000001010100;
reg [32-1:0] bias_reg_424 = 32'b00000000000000000000001010100000;
reg [32-1:0] bias_reg_425 = 32'b11111111111111111111111101110101;
reg [32-1:0] bias_reg_426 = 32'b11111111111111111111111110001011;
reg [32-1:0] bias_reg_427 = 32'b11111111111111111111111101101001;
reg [32-1:0] bias_reg_428 = 32'b11111111111111111111111111110110;
reg [32-1:0] bias_reg_429 = 32'b11111111111111111111111100001101;
reg [32-1:0] bias_reg_430 = 32'b11111111111111111111111110111000;
reg [32-1:0] bias_reg_431 = 32'b00000000000000000000000001111100;
reg [32-1:0] bias_reg_432 = 32'b00000000000000000000000001111111;
reg [32-1:0] bias_reg_433 = 32'b00000000000000000000000010001000;
reg [32-1:0] bias_reg_434 = 32'b11111111111111111111111110110011;
reg [32-1:0] bias_reg_435 = 32'b00000000000000000000000001000011;
reg [32-1:0] bias_reg_436 = 32'b00000000000000000000000011011101;
reg [32-1:0] bias_reg_437 = 32'b11111111111111111111111100110011;
reg [32-1:0] bias_reg_438 = 32'b11111111111111111111111101010101;
reg [32-1:0] bias_reg_439 = 32'b11111111111111111111111110001111;
reg [32-1:0] bias_reg_440 = 32'b00000000000000000000000010000011;
reg [32-1:0] bias_reg_441 = 32'b00000000000000000000000010101011;
reg [32-1:0] bias_reg_442 = 32'b11111111111111111111111111001010;
reg [32-1:0] bias_reg_443 = 32'b00000000000000000000001010101001;
reg [32-1:0] bias_reg_444 = 32'b00000000000000000000000000000100;
reg [32-1:0] bias_reg_445 = 32'b00000000000000000000000101011100;
reg [32-1:0] bias_reg_446 = 32'b00000000000000000000001011110110;
reg [32-1:0] bias_reg_447 = 32'b11111111111111111111111010011100;
reg [32-1:0] bias_reg_448 = 32'b00000000000000000000000100011000;
reg [32-1:0] bias_reg_449 = 32'b11111111111111111111111111011011;
reg [32-1:0] bias_reg_450 = 32'b00000000000000000000000011100111;
reg [32-1:0] bias_reg_451 = 32'b11111111111111111111111111100100;
reg [32-1:0] bias_reg_452 = 32'b00000000000000000000000000100110;
reg [32-1:0] bias_reg_453 = 32'b00000000000000000000000101000100;
reg [32-1:0] bias_reg_454 = 32'b00000000000000000000001000001110;
reg [32-1:0] bias_reg_455 = 32'b00000000000000000000001010101011;
reg [32-1:0] bias_reg_456 = 32'b00000000000000000000000001110000;
reg [32-1:0] bias_reg_457 = 32'b00000000000000000000000101011111;
reg [32-1:0] bias_reg_458 = 32'b00000000000000000000000111111010;
reg [32-1:0] bias_reg_459 = 32'b00000000000000000000000001011000;
reg [32-1:0] bias_reg_460 = 32'b00000000000000000000000010010011;
reg [32-1:0] bias_reg_461 = 32'b11111111111111111111111011111110;
reg [32-1:0] bias_reg_462 = 32'b11111111111111111111111101100001;
reg [32-1:0] bias_reg_463 = 32'b11111111111111111111111100110011;
reg [32-1:0] bias_reg_464 = 32'b00000000000000000000001000011010;
reg [32-1:0] bias_reg_465 = 32'b11111111111111111111111100101101;
reg [32-1:0] bias_reg_466 = 32'b11111111111111111111111101101111;
reg [32-1:0] bias_reg_467 = 32'b00000000000000000000000000100111;
reg [32-1:0] bias_reg_468 = 32'b00000000000000000000000010101010;
reg [32-1:0] bias_reg_469 = 32'b11111111111111111111111000010001;
reg [32-1:0] bias_reg_470 = 32'b11111111111111111111111011101000;
reg [32-1:0] bias_reg_471 = 32'b11111111111111111111111101101100;
reg [32-1:0] bias_reg_472 = 32'b11111111111111111111111011011100;
reg [32-1:0] bias_reg_473 = 32'b11111111111111111111111010010100;
reg [32-1:0] bias_reg_474 = 32'b00000000000000000000001000001001;
reg [32-1:0] bias_reg_475 = 32'b11111111111111111111111110100110;
reg [32-1:0] bias_reg_476 = 32'b11111111111111111111111111010001;
reg [32-1:0] bias_reg_477 = 32'b00000000000000000000000000101000;
reg [32-1:0] bias_reg_478 = 32'b00000000000000000000001001001000;
reg [32-1:0] bias_reg_479 = 32'b11111111111111111111111100011010;
reg [32-1:0] bias_reg_480 = 32'b00000000000000000000001000000101;
reg [32-1:0] bias_reg_481 = 32'b00000000000000000000000011010000;
reg [32-1:0] bias_reg_482 = 32'b11111111111111111111111010000111;
reg [32-1:0] bias_reg_483 = 32'b11111111111111111111111101001111;
reg [32-1:0] bias_reg_484 = 32'b11111111111111111111111110111011;
reg [32-1:0] bias_reg_485 = 32'b11111111111111111111111110000010;
reg [32-1:0] bias_reg_486 = 32'b11111111111111111111111110110101;
reg [32-1:0] bias_reg_487 = 32'b00000000000000000000000001111100;
reg [32-1:0] bias_reg_488 = 32'b00000000000000000000000000101000;
reg [32-1:0] bias_reg_489 = 32'b00000000000000000000001001101110;
reg [32-1:0] bias_reg_490 = 32'b11111111111111111111111110011001;
reg [32-1:0] bias_reg_491 = 32'b00000000000000000000000010111110;
reg [32-1:0] bias_reg_492 = 32'b00000000000000000000000100011100;
reg [32-1:0] bias_reg_493 = 32'b00000000000000000000000001011100;
reg [32-1:0] bias_reg_494 = 32'b11111111111111111111111001001111;
reg [32-1:0] bias_reg_495 = 32'b00000000000000000000001001110000;
reg [32-1:0] bias_reg_496 = 32'b00000000000000000000000000111110;
reg [32-1:0] bias_reg_497 = 32'b11111111111111111111110111010111;
reg [32-1:0] bias_reg_498 = 32'b00000000000000000000000001000010;
reg [32-1:0] bias_reg_499 = 32'b11111111111111111111111100011011;
reg [32-1:0] bias_reg_500 = 32'b00000000000000000000001000101110;
reg [32-1:0] bias_reg_501 = 32'b11111111111111111111111011000001;
reg [32-1:0] bias_reg_502 = 32'b11111111111111111111111111111111;
reg [32-1:0] bias_reg_503 = 32'b11111111111111111111111010101001;
reg [32-1:0] bias_reg_504 = 32'b11111111111111111111111101011011;
reg [32-1:0] bias_reg_505 = 32'b11111111111111111111111110101000;
reg [32-1:0] bias_reg_506 = 32'b00000000000000000000000001101111;
reg [32-1:0] bias_reg_507 = 32'b11111111111111111111111010000111;
reg [32-1:0] bias_reg_508 = 32'b00000000000000000000000010001011;
reg [32-1:0] bias_reg_509 = 32'b00000000000000000000000101011101;
reg [32-1:0] bias_reg_510 = 32'b00000000000000000000000001001001;
reg [32-1:0] bias_reg_511 = 32'b00000000000000000000000100101011;
assign bias_mem[0] = bias_reg_0;
assign bias_mem[1] = bias_reg_1;
assign bias_mem[2] = bias_reg_2;
assign bias_mem[3] = bias_reg_3;
assign bias_mem[4] = bias_reg_4;
assign bias_mem[5] = bias_reg_5;
assign bias_mem[6] = bias_reg_6;
assign bias_mem[7] = bias_reg_7;
assign bias_mem[8] = bias_reg_8;
assign bias_mem[9] = bias_reg_9;
assign bias_mem[10] = bias_reg_10;
assign bias_mem[11] = bias_reg_11;
assign bias_mem[12] = bias_reg_12;
assign bias_mem[13] = bias_reg_13;
assign bias_mem[14] = bias_reg_14;
assign bias_mem[15] = bias_reg_15;
assign bias_mem[16] = bias_reg_16;
assign bias_mem[17] = bias_reg_17;
assign bias_mem[18] = bias_reg_18;
assign bias_mem[19] = bias_reg_19;
assign bias_mem[20] = bias_reg_20;
assign bias_mem[21] = bias_reg_21;
assign bias_mem[22] = bias_reg_22;
assign bias_mem[23] = bias_reg_23;
assign bias_mem[24] = bias_reg_24;
assign bias_mem[25] = bias_reg_25;
assign bias_mem[26] = bias_reg_26;
assign bias_mem[27] = bias_reg_27;
assign bias_mem[28] = bias_reg_28;
assign bias_mem[29] = bias_reg_29;
assign bias_mem[30] = bias_reg_30;
assign bias_mem[31] = bias_reg_31;
assign bias_mem[32] = bias_reg_32;
assign bias_mem[33] = bias_reg_33;
assign bias_mem[34] = bias_reg_34;
assign bias_mem[35] = bias_reg_35;
assign bias_mem[36] = bias_reg_36;
assign bias_mem[37] = bias_reg_37;
assign bias_mem[38] = bias_reg_38;
assign bias_mem[39] = bias_reg_39;
assign bias_mem[40] = bias_reg_40;
assign bias_mem[41] = bias_reg_41;
assign bias_mem[42] = bias_reg_42;
assign bias_mem[43] = bias_reg_43;
assign bias_mem[44] = bias_reg_44;
assign bias_mem[45] = bias_reg_45;
assign bias_mem[46] = bias_reg_46;
assign bias_mem[47] = bias_reg_47;
assign bias_mem[48] = bias_reg_48;
assign bias_mem[49] = bias_reg_49;
assign bias_mem[50] = bias_reg_50;
assign bias_mem[51] = bias_reg_51;
assign bias_mem[52] = bias_reg_52;
assign bias_mem[53] = bias_reg_53;
assign bias_mem[54] = bias_reg_54;
assign bias_mem[55] = bias_reg_55;
assign bias_mem[56] = bias_reg_56;
assign bias_mem[57] = bias_reg_57;
assign bias_mem[58] = bias_reg_58;
assign bias_mem[59] = bias_reg_59;
assign bias_mem[60] = bias_reg_60;
assign bias_mem[61] = bias_reg_61;
assign bias_mem[62] = bias_reg_62;
assign bias_mem[63] = bias_reg_63;
assign bias_mem[64] = bias_reg_64;
assign bias_mem[65] = bias_reg_65;
assign bias_mem[66] = bias_reg_66;
assign bias_mem[67] = bias_reg_67;
assign bias_mem[68] = bias_reg_68;
assign bias_mem[69] = bias_reg_69;
assign bias_mem[70] = bias_reg_70;
assign bias_mem[71] = bias_reg_71;
assign bias_mem[72] = bias_reg_72;
assign bias_mem[73] = bias_reg_73;
assign bias_mem[74] = bias_reg_74;
assign bias_mem[75] = bias_reg_75;
assign bias_mem[76] = bias_reg_76;
assign bias_mem[77] = bias_reg_77;
assign bias_mem[78] = bias_reg_78;
assign bias_mem[79] = bias_reg_79;
assign bias_mem[80] = bias_reg_80;
assign bias_mem[81] = bias_reg_81;
assign bias_mem[82] = bias_reg_82;
assign bias_mem[83] = bias_reg_83;
assign bias_mem[84] = bias_reg_84;
assign bias_mem[85] = bias_reg_85;
assign bias_mem[86] = bias_reg_86;
assign bias_mem[87] = bias_reg_87;
assign bias_mem[88] = bias_reg_88;
assign bias_mem[89] = bias_reg_89;
assign bias_mem[90] = bias_reg_90;
assign bias_mem[91] = bias_reg_91;
assign bias_mem[92] = bias_reg_92;
assign bias_mem[93] = bias_reg_93;
assign bias_mem[94] = bias_reg_94;
assign bias_mem[95] = bias_reg_95;
assign bias_mem[96] = bias_reg_96;
assign bias_mem[97] = bias_reg_97;
assign bias_mem[98] = bias_reg_98;
assign bias_mem[99] = bias_reg_99;
assign bias_mem[100] = bias_reg_100;
assign bias_mem[101] = bias_reg_101;
assign bias_mem[102] = bias_reg_102;
assign bias_mem[103] = bias_reg_103;
assign bias_mem[104] = bias_reg_104;
assign bias_mem[105] = bias_reg_105;
assign bias_mem[106] = bias_reg_106;
assign bias_mem[107] = bias_reg_107;
assign bias_mem[108] = bias_reg_108;
assign bias_mem[109] = bias_reg_109;
assign bias_mem[110] = bias_reg_110;
assign bias_mem[111] = bias_reg_111;
assign bias_mem[112] = bias_reg_112;
assign bias_mem[113] = bias_reg_113;
assign bias_mem[114] = bias_reg_114;
assign bias_mem[115] = bias_reg_115;
assign bias_mem[116] = bias_reg_116;
assign bias_mem[117] = bias_reg_117;
assign bias_mem[118] = bias_reg_118;
assign bias_mem[119] = bias_reg_119;
assign bias_mem[120] = bias_reg_120;
assign bias_mem[121] = bias_reg_121;
assign bias_mem[122] = bias_reg_122;
assign bias_mem[123] = bias_reg_123;
assign bias_mem[124] = bias_reg_124;
assign bias_mem[125] = bias_reg_125;
assign bias_mem[126] = bias_reg_126;
assign bias_mem[127] = bias_reg_127;
assign bias_mem[128] = bias_reg_128;
assign bias_mem[129] = bias_reg_129;
assign bias_mem[130] = bias_reg_130;
assign bias_mem[131] = bias_reg_131;
assign bias_mem[132] = bias_reg_132;
assign bias_mem[133] = bias_reg_133;
assign bias_mem[134] = bias_reg_134;
assign bias_mem[135] = bias_reg_135;
assign bias_mem[136] = bias_reg_136;
assign bias_mem[137] = bias_reg_137;
assign bias_mem[138] = bias_reg_138;
assign bias_mem[139] = bias_reg_139;
assign bias_mem[140] = bias_reg_140;
assign bias_mem[141] = bias_reg_141;
assign bias_mem[142] = bias_reg_142;
assign bias_mem[143] = bias_reg_143;
assign bias_mem[144] = bias_reg_144;
assign bias_mem[145] = bias_reg_145;
assign bias_mem[146] = bias_reg_146;
assign bias_mem[147] = bias_reg_147;
assign bias_mem[148] = bias_reg_148;
assign bias_mem[149] = bias_reg_149;
assign bias_mem[150] = bias_reg_150;
assign bias_mem[151] = bias_reg_151;
assign bias_mem[152] = bias_reg_152;
assign bias_mem[153] = bias_reg_153;
assign bias_mem[154] = bias_reg_154;
assign bias_mem[155] = bias_reg_155;
assign bias_mem[156] = bias_reg_156;
assign bias_mem[157] = bias_reg_157;
assign bias_mem[158] = bias_reg_158;
assign bias_mem[159] = bias_reg_159;
assign bias_mem[160] = bias_reg_160;
assign bias_mem[161] = bias_reg_161;
assign bias_mem[162] = bias_reg_162;
assign bias_mem[163] = bias_reg_163;
assign bias_mem[164] = bias_reg_164;
assign bias_mem[165] = bias_reg_165;
assign bias_mem[166] = bias_reg_166;
assign bias_mem[167] = bias_reg_167;
assign bias_mem[168] = bias_reg_168;
assign bias_mem[169] = bias_reg_169;
assign bias_mem[170] = bias_reg_170;
assign bias_mem[171] = bias_reg_171;
assign bias_mem[172] = bias_reg_172;
assign bias_mem[173] = bias_reg_173;
assign bias_mem[174] = bias_reg_174;
assign bias_mem[175] = bias_reg_175;
assign bias_mem[176] = bias_reg_176;
assign bias_mem[177] = bias_reg_177;
assign bias_mem[178] = bias_reg_178;
assign bias_mem[179] = bias_reg_179;
assign bias_mem[180] = bias_reg_180;
assign bias_mem[181] = bias_reg_181;
assign bias_mem[182] = bias_reg_182;
assign bias_mem[183] = bias_reg_183;
assign bias_mem[184] = bias_reg_184;
assign bias_mem[185] = bias_reg_185;
assign bias_mem[186] = bias_reg_186;
assign bias_mem[187] = bias_reg_187;
assign bias_mem[188] = bias_reg_188;
assign bias_mem[189] = bias_reg_189;
assign bias_mem[190] = bias_reg_190;
assign bias_mem[191] = bias_reg_191;
assign bias_mem[192] = bias_reg_192;
assign bias_mem[193] = bias_reg_193;
assign bias_mem[194] = bias_reg_194;
assign bias_mem[195] = bias_reg_195;
assign bias_mem[196] = bias_reg_196;
assign bias_mem[197] = bias_reg_197;
assign bias_mem[198] = bias_reg_198;
assign bias_mem[199] = bias_reg_199;
assign bias_mem[200] = bias_reg_200;
assign bias_mem[201] = bias_reg_201;
assign bias_mem[202] = bias_reg_202;
assign bias_mem[203] = bias_reg_203;
assign bias_mem[204] = bias_reg_204;
assign bias_mem[205] = bias_reg_205;
assign bias_mem[206] = bias_reg_206;
assign bias_mem[207] = bias_reg_207;
assign bias_mem[208] = bias_reg_208;
assign bias_mem[209] = bias_reg_209;
assign bias_mem[210] = bias_reg_210;
assign bias_mem[211] = bias_reg_211;
assign bias_mem[212] = bias_reg_212;
assign bias_mem[213] = bias_reg_213;
assign bias_mem[214] = bias_reg_214;
assign bias_mem[215] = bias_reg_215;
assign bias_mem[216] = bias_reg_216;
assign bias_mem[217] = bias_reg_217;
assign bias_mem[218] = bias_reg_218;
assign bias_mem[219] = bias_reg_219;
assign bias_mem[220] = bias_reg_220;
assign bias_mem[221] = bias_reg_221;
assign bias_mem[222] = bias_reg_222;
assign bias_mem[223] = bias_reg_223;
assign bias_mem[224] = bias_reg_224;
assign bias_mem[225] = bias_reg_225;
assign bias_mem[226] = bias_reg_226;
assign bias_mem[227] = bias_reg_227;
assign bias_mem[228] = bias_reg_228;
assign bias_mem[229] = bias_reg_229;
assign bias_mem[230] = bias_reg_230;
assign bias_mem[231] = bias_reg_231;
assign bias_mem[232] = bias_reg_232;
assign bias_mem[233] = bias_reg_233;
assign bias_mem[234] = bias_reg_234;
assign bias_mem[235] = bias_reg_235;
assign bias_mem[236] = bias_reg_236;
assign bias_mem[237] = bias_reg_237;
assign bias_mem[238] = bias_reg_238;
assign bias_mem[239] = bias_reg_239;
assign bias_mem[240] = bias_reg_240;
assign bias_mem[241] = bias_reg_241;
assign bias_mem[242] = bias_reg_242;
assign bias_mem[243] = bias_reg_243;
assign bias_mem[244] = bias_reg_244;
assign bias_mem[245] = bias_reg_245;
assign bias_mem[246] = bias_reg_246;
assign bias_mem[247] = bias_reg_247;
assign bias_mem[248] = bias_reg_248;
assign bias_mem[249] = bias_reg_249;
assign bias_mem[250] = bias_reg_250;
assign bias_mem[251] = bias_reg_251;
assign bias_mem[252] = bias_reg_252;
assign bias_mem[253] = bias_reg_253;
assign bias_mem[254] = bias_reg_254;
assign bias_mem[255] = bias_reg_255;
assign bias_mem[256] = bias_reg_256;
assign bias_mem[257] = bias_reg_257;
assign bias_mem[258] = bias_reg_258;
assign bias_mem[259] = bias_reg_259;
assign bias_mem[260] = bias_reg_260;
assign bias_mem[261] = bias_reg_261;
assign bias_mem[262] = bias_reg_262;
assign bias_mem[263] = bias_reg_263;
assign bias_mem[264] = bias_reg_264;
assign bias_mem[265] = bias_reg_265;
assign bias_mem[266] = bias_reg_266;
assign bias_mem[267] = bias_reg_267;
assign bias_mem[268] = bias_reg_268;
assign bias_mem[269] = bias_reg_269;
assign bias_mem[270] = bias_reg_270;
assign bias_mem[271] = bias_reg_271;
assign bias_mem[272] = bias_reg_272;
assign bias_mem[273] = bias_reg_273;
assign bias_mem[274] = bias_reg_274;
assign bias_mem[275] = bias_reg_275;
assign bias_mem[276] = bias_reg_276;
assign bias_mem[277] = bias_reg_277;
assign bias_mem[278] = bias_reg_278;
assign bias_mem[279] = bias_reg_279;
assign bias_mem[280] = bias_reg_280;
assign bias_mem[281] = bias_reg_281;
assign bias_mem[282] = bias_reg_282;
assign bias_mem[283] = bias_reg_283;
assign bias_mem[284] = bias_reg_284;
assign bias_mem[285] = bias_reg_285;
assign bias_mem[286] = bias_reg_286;
assign bias_mem[287] = bias_reg_287;
assign bias_mem[288] = bias_reg_288;
assign bias_mem[289] = bias_reg_289;
assign bias_mem[290] = bias_reg_290;
assign bias_mem[291] = bias_reg_291;
assign bias_mem[292] = bias_reg_292;
assign bias_mem[293] = bias_reg_293;
assign bias_mem[294] = bias_reg_294;
assign bias_mem[295] = bias_reg_295;
assign bias_mem[296] = bias_reg_296;
assign bias_mem[297] = bias_reg_297;
assign bias_mem[298] = bias_reg_298;
assign bias_mem[299] = bias_reg_299;
assign bias_mem[300] = bias_reg_300;
assign bias_mem[301] = bias_reg_301;
assign bias_mem[302] = bias_reg_302;
assign bias_mem[303] = bias_reg_303;
assign bias_mem[304] = bias_reg_304;
assign bias_mem[305] = bias_reg_305;
assign bias_mem[306] = bias_reg_306;
assign bias_mem[307] = bias_reg_307;
assign bias_mem[308] = bias_reg_308;
assign bias_mem[309] = bias_reg_309;
assign bias_mem[310] = bias_reg_310;
assign bias_mem[311] = bias_reg_311;
assign bias_mem[312] = bias_reg_312;
assign bias_mem[313] = bias_reg_313;
assign bias_mem[314] = bias_reg_314;
assign bias_mem[315] = bias_reg_315;
assign bias_mem[316] = bias_reg_316;
assign bias_mem[317] = bias_reg_317;
assign bias_mem[318] = bias_reg_318;
assign bias_mem[319] = bias_reg_319;
assign bias_mem[320] = bias_reg_320;
assign bias_mem[321] = bias_reg_321;
assign bias_mem[322] = bias_reg_322;
assign bias_mem[323] = bias_reg_323;
assign bias_mem[324] = bias_reg_324;
assign bias_mem[325] = bias_reg_325;
assign bias_mem[326] = bias_reg_326;
assign bias_mem[327] = bias_reg_327;
assign bias_mem[328] = bias_reg_328;
assign bias_mem[329] = bias_reg_329;
assign bias_mem[330] = bias_reg_330;
assign bias_mem[331] = bias_reg_331;
assign bias_mem[332] = bias_reg_332;
assign bias_mem[333] = bias_reg_333;
assign bias_mem[334] = bias_reg_334;
assign bias_mem[335] = bias_reg_335;
assign bias_mem[336] = bias_reg_336;
assign bias_mem[337] = bias_reg_337;
assign bias_mem[338] = bias_reg_338;
assign bias_mem[339] = bias_reg_339;
assign bias_mem[340] = bias_reg_340;
assign bias_mem[341] = bias_reg_341;
assign bias_mem[342] = bias_reg_342;
assign bias_mem[343] = bias_reg_343;
assign bias_mem[344] = bias_reg_344;
assign bias_mem[345] = bias_reg_345;
assign bias_mem[346] = bias_reg_346;
assign bias_mem[347] = bias_reg_347;
assign bias_mem[348] = bias_reg_348;
assign bias_mem[349] = bias_reg_349;
assign bias_mem[350] = bias_reg_350;
assign bias_mem[351] = bias_reg_351;
assign bias_mem[352] = bias_reg_352;
assign bias_mem[353] = bias_reg_353;
assign bias_mem[354] = bias_reg_354;
assign bias_mem[355] = bias_reg_355;
assign bias_mem[356] = bias_reg_356;
assign bias_mem[357] = bias_reg_357;
assign bias_mem[358] = bias_reg_358;
assign bias_mem[359] = bias_reg_359;
assign bias_mem[360] = bias_reg_360;
assign bias_mem[361] = bias_reg_361;
assign bias_mem[362] = bias_reg_362;
assign bias_mem[363] = bias_reg_363;
assign bias_mem[364] = bias_reg_364;
assign bias_mem[365] = bias_reg_365;
assign bias_mem[366] = bias_reg_366;
assign bias_mem[367] = bias_reg_367;
assign bias_mem[368] = bias_reg_368;
assign bias_mem[369] = bias_reg_369;
assign bias_mem[370] = bias_reg_370;
assign bias_mem[371] = bias_reg_371;
assign bias_mem[372] = bias_reg_372;
assign bias_mem[373] = bias_reg_373;
assign bias_mem[374] = bias_reg_374;
assign bias_mem[375] = bias_reg_375;
assign bias_mem[376] = bias_reg_376;
assign bias_mem[377] = bias_reg_377;
assign bias_mem[378] = bias_reg_378;
assign bias_mem[379] = bias_reg_379;
assign bias_mem[380] = bias_reg_380;
assign bias_mem[381] = bias_reg_381;
assign bias_mem[382] = bias_reg_382;
assign bias_mem[383] = bias_reg_383;
assign bias_mem[384] = bias_reg_384;
assign bias_mem[385] = bias_reg_385;
assign bias_mem[386] = bias_reg_386;
assign bias_mem[387] = bias_reg_387;
assign bias_mem[388] = bias_reg_388;
assign bias_mem[389] = bias_reg_389;
assign bias_mem[390] = bias_reg_390;
assign bias_mem[391] = bias_reg_391;
assign bias_mem[392] = bias_reg_392;
assign bias_mem[393] = bias_reg_393;
assign bias_mem[394] = bias_reg_394;
assign bias_mem[395] = bias_reg_395;
assign bias_mem[396] = bias_reg_396;
assign bias_mem[397] = bias_reg_397;
assign bias_mem[398] = bias_reg_398;
assign bias_mem[399] = bias_reg_399;
assign bias_mem[400] = bias_reg_400;
assign bias_mem[401] = bias_reg_401;
assign bias_mem[402] = bias_reg_402;
assign bias_mem[403] = bias_reg_403;
assign bias_mem[404] = bias_reg_404;
assign bias_mem[405] = bias_reg_405;
assign bias_mem[406] = bias_reg_406;
assign bias_mem[407] = bias_reg_407;
assign bias_mem[408] = bias_reg_408;
assign bias_mem[409] = bias_reg_409;
assign bias_mem[410] = bias_reg_410;
assign bias_mem[411] = bias_reg_411;
assign bias_mem[412] = bias_reg_412;
assign bias_mem[413] = bias_reg_413;
assign bias_mem[414] = bias_reg_414;
assign bias_mem[415] = bias_reg_415;
assign bias_mem[416] = bias_reg_416;
assign bias_mem[417] = bias_reg_417;
assign bias_mem[418] = bias_reg_418;
assign bias_mem[419] = bias_reg_419;
assign bias_mem[420] = bias_reg_420;
assign bias_mem[421] = bias_reg_421;
assign bias_mem[422] = bias_reg_422;
assign bias_mem[423] = bias_reg_423;
assign bias_mem[424] = bias_reg_424;
assign bias_mem[425] = bias_reg_425;
assign bias_mem[426] = bias_reg_426;
assign bias_mem[427] = bias_reg_427;
assign bias_mem[428] = bias_reg_428;
assign bias_mem[429] = bias_reg_429;
assign bias_mem[430] = bias_reg_430;
assign bias_mem[431] = bias_reg_431;
assign bias_mem[432] = bias_reg_432;
assign bias_mem[433] = bias_reg_433;
assign bias_mem[434] = bias_reg_434;
assign bias_mem[435] = bias_reg_435;
assign bias_mem[436] = bias_reg_436;
assign bias_mem[437] = bias_reg_437;
assign bias_mem[438] = bias_reg_438;
assign bias_mem[439] = bias_reg_439;
assign bias_mem[440] = bias_reg_440;
assign bias_mem[441] = bias_reg_441;
assign bias_mem[442] = bias_reg_442;
assign bias_mem[443] = bias_reg_443;
assign bias_mem[444] = bias_reg_444;
assign bias_mem[445] = bias_reg_445;
assign bias_mem[446] = bias_reg_446;
assign bias_mem[447] = bias_reg_447;
assign bias_mem[448] = bias_reg_448;
assign bias_mem[449] = bias_reg_449;
assign bias_mem[450] = bias_reg_450;
assign bias_mem[451] = bias_reg_451;
assign bias_mem[452] = bias_reg_452;
assign bias_mem[453] = bias_reg_453;
assign bias_mem[454] = bias_reg_454;
assign bias_mem[455] = bias_reg_455;
assign bias_mem[456] = bias_reg_456;
assign bias_mem[457] = bias_reg_457;
assign bias_mem[458] = bias_reg_458;
assign bias_mem[459] = bias_reg_459;
assign bias_mem[460] = bias_reg_460;
assign bias_mem[461] = bias_reg_461;
assign bias_mem[462] = bias_reg_462;
assign bias_mem[463] = bias_reg_463;
assign bias_mem[464] = bias_reg_464;
assign bias_mem[465] = bias_reg_465;
assign bias_mem[466] = bias_reg_466;
assign bias_mem[467] = bias_reg_467;
assign bias_mem[468] = bias_reg_468;
assign bias_mem[469] = bias_reg_469;
assign bias_mem[470] = bias_reg_470;
assign bias_mem[471] = bias_reg_471;
assign bias_mem[472] = bias_reg_472;
assign bias_mem[473] = bias_reg_473;
assign bias_mem[474] = bias_reg_474;
assign bias_mem[475] = bias_reg_475;
assign bias_mem[476] = bias_reg_476;
assign bias_mem[477] = bias_reg_477;
assign bias_mem[478] = bias_reg_478;
assign bias_mem[479] = bias_reg_479;
assign bias_mem[480] = bias_reg_480;
assign bias_mem[481] = bias_reg_481;
assign bias_mem[482] = bias_reg_482;
assign bias_mem[483] = bias_reg_483;
assign bias_mem[484] = bias_reg_484;
assign bias_mem[485] = bias_reg_485;
assign bias_mem[486] = bias_reg_486;
assign bias_mem[487] = bias_reg_487;
assign bias_mem[488] = bias_reg_488;
assign bias_mem[489] = bias_reg_489;
assign bias_mem[490] = bias_reg_490;
assign bias_mem[491] = bias_reg_491;
assign bias_mem[492] = bias_reg_492;
assign bias_mem[493] = bias_reg_493;
assign bias_mem[494] = bias_reg_494;
assign bias_mem[495] = bias_reg_495;
assign bias_mem[496] = bias_reg_496;
assign bias_mem[497] = bias_reg_497;
assign bias_mem[498] = bias_reg_498;
assign bias_mem[499] = bias_reg_499;
assign bias_mem[500] = bias_reg_500;
assign bias_mem[501] = bias_reg_501;
assign bias_mem[502] = bias_reg_502;
assign bias_mem[503] = bias_reg_503;
assign bias_mem[504] = bias_reg_504;
assign bias_mem[505] = bias_reg_505;
assign bias_mem[506] = bias_reg_506;
assign bias_mem[507] = bias_reg_507;
assign bias_mem[508] = bias_reg_508;
assign bias_mem[509] = bias_reg_509;
assign bias_mem[510] = bias_reg_510;
assign bias_mem[511] = bias_reg_511;
endmodule
