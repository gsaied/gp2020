
	/* verilator lint_off COMBDLY */
	module rom_fire3_squeeze #(
	parameter WIDTH=16,
	parameter KERNEL=1,
	parameter ADDR=7,
	parameter NUM=16)
	(
		input [ADDR-1:0] address ,
		//input clk,
		output [WIDTH-1:0] rom_out [0:NUM-1]
	);	
	

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_1 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_2 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_3 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_4 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_5 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_6 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_7 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_8 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_9 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_10 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_11 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_12 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_13 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_14 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_15 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_16 [0:2**ADDR-1] ;
initial  begin
$readmemb("fire3_squeeze/file_fire3_squeeze_1.mem",rom_1,0,2**ADDR-1);
$readmemb("fire3_squeeze/file_fire3_squeeze_2.mem",rom_2,0,2**ADDR-1);
$readmemb("fire3_squeeze/file_fire3_squeeze_3.mem",rom_3,0,2**ADDR-1);
$readmemb("fire3_squeeze/file_fire3_squeeze_4.mem",rom_4,0,2**ADDR-1);
$readmemb("fire3_squeeze/file_fire3_squeeze_5.mem",rom_5,0,2**ADDR-1);
$readmemb("fire3_squeeze/file_fire3_squeeze_6.mem",rom_6,0,2**ADDR-1);
$readmemb("fire3_squeeze/file_fire3_squeeze_7.mem",rom_7,0,2**ADDR-1);
$readmemb("fire3_squeeze/file_fire3_squeeze_8.mem",rom_8,0,2**ADDR-1);
$readmemb("fire3_squeeze/file_fire3_squeeze_9.mem",rom_9,0,2**ADDR-1);
$readmemb("fire3_squeeze/file_fire3_squeeze_10.mem",rom_10,0,2**ADDR-1);
$readmemb("fire3_squeeze/file_fire3_squeeze_11.mem",rom_11,0,2**ADDR-1);
$readmemb("fire3_squeeze/file_fire3_squeeze_12.mem",rom_12,0,2**ADDR-1);
$readmemb("fire3_squeeze/file_fire3_squeeze_13.mem",rom_13,0,2**ADDR-1);
$readmemb("fire3_squeeze/file_fire3_squeeze_14.mem",rom_14,0,2**ADDR-1);
$readmemb("fire3_squeeze/file_fire3_squeeze_15.mem",rom_15,0,2**ADDR-1);
$readmemb("fire3_squeeze/file_fire3_squeeze_16.mem",rom_16,0,2**ADDR-1);
end
assign rom_out[0] = rom_1[address] ;
assign rom_out[1] = rom_2[address] ;
assign rom_out[2] = rom_3[address] ;
assign rom_out[3] = rom_4[address] ;
assign rom_out[4] = rom_5[address] ;
assign rom_out[5] = rom_6[address] ;
assign rom_out[6] = rom_7[address] ;
assign rom_out[7] = rom_8[address] ;
assign rom_out[8] = rom_9[address] ;
assign rom_out[9] = rom_10[address] ;
assign rom_out[10] = rom_11[address] ;
assign rom_out[11] = rom_12[address] ;
assign rom_out[12] = rom_13[address] ;
assign rom_out[13] = rom_14[address] ;
assign rom_out[14] = rom_15[address] ;
assign rom_out[15] = rom_16[address] ;
endmodule
