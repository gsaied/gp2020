module rom #(
	parameter WIDHT=16,
	parameter NUM=4
)
(
	input clk,
	input address,
	output reg [WIDTH-1:0] kernel
);


endmodule
