
module biasing_fire4_squeeze (
	output [32-1:0] bias_mem [0:32-1]
);

reg [32-1:0] bias_reg_0 = 32'b00000000000000000000000101100000;
reg [32-1:0] bias_reg_1 = 32'b00000000000000000000010000100000;
reg [32-1:0] bias_reg_2 = 32'b00000000000000000000000001100000;
reg [32-1:0] bias_reg_3 = 32'b00000000000000000000000010111010;
reg [32-1:0] bias_reg_4 = 32'b00000000000000000000000100111011;
reg [32-1:0] bias_reg_5 = 32'b11111111111111111111111011111001;
reg [32-1:0] bias_reg_6 = 32'b11111111111111111111111001110100;
reg [32-1:0] bias_reg_7 = 32'b11111111111111111111111100111101;
reg [32-1:0] bias_reg_8 = 32'b11111111111111111111111111001100;
reg [32-1:0] bias_reg_9 = 32'b11111111111111111111111101101011;
reg [32-1:0] bias_reg_10 = 32'b11111111111111111111111110010111;
reg [32-1:0] bias_reg_11 = 32'b00000000000000000000000001011001;
reg [32-1:0] bias_reg_12 = 32'b00000000000000000000000001011110;
reg [32-1:0] bias_reg_13 = 32'b00000000000000000000000011111101;
reg [32-1:0] bias_reg_14 = 32'b00000000000000000000000011011101;
reg [32-1:0] bias_reg_15 = 32'b00000000000000000000000000011001;
reg [32-1:0] bias_reg_16 = 32'b00000000000000000000001011000000;
reg [32-1:0] bias_reg_17 = 32'b00000000000000000000001000101101;
reg [32-1:0] bias_reg_18 = 32'b00000000000000000000000110011011;
reg [32-1:0] bias_reg_19 = 32'b00000000000000000000000000011111;
reg [32-1:0] bias_reg_20 = 32'b11111111111111111111111100001111;
reg [32-1:0] bias_reg_21 = 32'b00000000000000000000000000110010;
reg [32-1:0] bias_reg_22 = 32'b11111111111111111111110111100011;
reg [32-1:0] bias_reg_23 = 32'b00000000000000000000001001011101;
reg [32-1:0] bias_reg_24 = 32'b00000000000000000000000110100000;
reg [32-1:0] bias_reg_25 = 32'b00000000000000000000000000111101;
reg [32-1:0] bias_reg_26 = 32'b00000000000000000000000000000000;
reg [32-1:0] bias_reg_27 = 32'b00000000000000000000000111111110;
reg [32-1:0] bias_reg_28 = 32'b00000000000000000000000100001000;
reg [32-1:0] bias_reg_29 = 32'b11111111111111111111110101011110;
reg [32-1:0] bias_reg_30 = 32'b00000000000000000000000001100110;
reg [32-1:0] bias_reg_31 = 32'b11111111111111111111111010010110;
assign bias_mem[0] = bias_reg_0;
assign bias_mem[1] = bias_reg_1;
assign bias_mem[2] = bias_reg_2;
assign bias_mem[3] = bias_reg_3;
assign bias_mem[4] = bias_reg_4;
assign bias_mem[5] = bias_reg_5;
assign bias_mem[6] = bias_reg_6;
assign bias_mem[7] = bias_reg_7;
assign bias_mem[8] = bias_reg_8;
assign bias_mem[9] = bias_reg_9;
assign bias_mem[10] = bias_reg_10;
assign bias_mem[11] = bias_reg_11;
assign bias_mem[12] = bias_reg_12;
assign bias_mem[13] = bias_reg_13;
assign bias_mem[14] = bias_reg_14;
assign bias_mem[15] = bias_reg_15;
assign bias_mem[16] = bias_reg_16;
assign bias_mem[17] = bias_reg_17;
assign bias_mem[18] = bias_reg_18;
assign bias_mem[19] = bias_reg_19;
assign bias_mem[20] = bias_reg_20;
assign bias_mem[21] = bias_reg_21;
assign bias_mem[22] = bias_reg_22;
assign bias_mem[23] = bias_reg_23;
assign bias_mem[24] = bias_reg_24;
assign bias_mem[25] = bias_reg_25;
assign bias_mem[26] = bias_reg_26;
assign bias_mem[27] = bias_reg_27;
assign bias_mem[28] = bias_reg_28;
assign bias_mem[29] = bias_reg_29;
assign bias_mem[30] = bias_reg_30;
assign bias_mem[31] = bias_reg_31;
endmodule
