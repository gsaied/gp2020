
module biasing_fire4_expand3 (
	output [32-1:0] bias_mem [0:128-1]
);

reg [32-1:0] bias_reg_0 = 32'b11111111111111111111111111000011;
reg [32-1:0] bias_reg_1 = 32'b00000000000000000000000000010101;
reg [32-1:0] bias_reg_2 = 32'b11111111111111111111111111000100;
reg [32-1:0] bias_reg_3 = 32'b00000000000000000000000100001010;
reg [32-1:0] bias_reg_4 = 32'b00000000000000000000000010000111;
reg [32-1:0] bias_reg_5 = 32'b11111111111111111111111110000110;
reg [32-1:0] bias_reg_6 = 32'b00000000000000000000000001011001;
reg [32-1:0] bias_reg_7 = 32'b00000000000000000000000000100110;
reg [32-1:0] bias_reg_8 = 32'b11111111111111111111111111000011;
reg [32-1:0] bias_reg_9 = 32'b11111111111111111111111111110000;
reg [32-1:0] bias_reg_10 = 32'b11111111111111111111111111110101;
reg [32-1:0] bias_reg_11 = 32'b00000000000000000000000000011111;
reg [32-1:0] bias_reg_12 = 32'b11111111111111111111111111001000;
reg [32-1:0] bias_reg_13 = 32'b11111111111111111111111111010110;
reg [32-1:0] bias_reg_14 = 32'b00000000000000000000000010011000;
reg [32-1:0] bias_reg_15 = 32'b11111111111111111111111111111011;
reg [32-1:0] bias_reg_16 = 32'b00000000000000000000000100010111;
reg [32-1:0] bias_reg_17 = 32'b11111111111111111111111111101000;
reg [32-1:0] bias_reg_18 = 32'b00000000000000000000000000001100;
reg [32-1:0] bias_reg_19 = 32'b00000000000000000000000000000101;
reg [32-1:0] bias_reg_20 = 32'b00000000000000000000000011110011;
reg [32-1:0] bias_reg_21 = 32'b00000000000000000000000000010000;
reg [32-1:0] bias_reg_22 = 32'b11111111111111111111111111010100;
reg [32-1:0] bias_reg_23 = 32'b00000000000000000000000000000110;
reg [32-1:0] bias_reg_24 = 32'b11111111111111111111111111100011;
reg [32-1:0] bias_reg_25 = 32'b11111111111111111111111111010101;
reg [32-1:0] bias_reg_26 = 32'b11111111111111111111111111001011;
reg [32-1:0] bias_reg_27 = 32'b00000000000000000000000010010100;
reg [32-1:0] bias_reg_28 = 32'b11111111111111111111111111100010;
reg [32-1:0] bias_reg_29 = 32'b00000000000000000000000010101011;
reg [32-1:0] bias_reg_30 = 32'b11111111111111111111111111001011;
reg [32-1:0] bias_reg_31 = 32'b11111111111111111111111111111101;
reg [32-1:0] bias_reg_32 = 32'b11111111111111111111111111010000;
reg [32-1:0] bias_reg_33 = 32'b11111111111111111111111110100100;
reg [32-1:0] bias_reg_34 = 32'b11111111111111111111111111100101;
reg [32-1:0] bias_reg_35 = 32'b00000000000000000000000001011100;
reg [32-1:0] bias_reg_36 = 32'b11111111111111111111111111100001;
reg [32-1:0] bias_reg_37 = 32'b00000000000000000000000000111010;
reg [32-1:0] bias_reg_38 = 32'b00000000000000000000000001001101;
reg [32-1:0] bias_reg_39 = 32'b11111111111111111111111111101111;
reg [32-1:0] bias_reg_40 = 32'b00000000000000000000000000011110;
reg [32-1:0] bias_reg_41 = 32'b11111111111111111111111111011111;
reg [32-1:0] bias_reg_42 = 32'b11111111111111111111111111101111;
reg [32-1:0] bias_reg_43 = 32'b00000000000000000000000001010010;
reg [32-1:0] bias_reg_44 = 32'b11111111111111111111111111111100;
reg [32-1:0] bias_reg_45 = 32'b11111111111111111111111110111001;
reg [32-1:0] bias_reg_46 = 32'b00000000000000000000000000001010;
reg [32-1:0] bias_reg_47 = 32'b00000000000000000000000000000001;
reg [32-1:0] bias_reg_48 = 32'b11111111111111111111111111110111;
reg [32-1:0] bias_reg_49 = 32'b11111111111111111111111111000110;
reg [32-1:0] bias_reg_50 = 32'b11111111111111111111111111100111;
reg [32-1:0] bias_reg_51 = 32'b00000000000000000000000000000010;
reg [32-1:0] bias_reg_52 = 32'b00000000000000000000000000011101;
reg [32-1:0] bias_reg_53 = 32'b11111111111111111111111111010000;
reg [32-1:0] bias_reg_54 = 32'b00000000000000000000000000010101;
reg [32-1:0] bias_reg_55 = 32'b00000000000000000000000000000101;
reg [32-1:0] bias_reg_56 = 32'b11111111111111111111111110111100;
reg [32-1:0] bias_reg_57 = 32'b00000000000000000000000000000010;
reg [32-1:0] bias_reg_58 = 32'b00000000000000000000000000000010;
reg [32-1:0] bias_reg_59 = 32'b11111111111111111111111111100010;
reg [32-1:0] bias_reg_60 = 32'b11111111111111111111111111100011;
reg [32-1:0] bias_reg_61 = 32'b11111111111111111111111110110010;
reg [32-1:0] bias_reg_62 = 32'b11111111111111111111111111110101;
reg [32-1:0] bias_reg_63 = 32'b00000000000000000000000011110001;
reg [32-1:0] bias_reg_64 = 32'b11111111111111111111111111100101;
reg [32-1:0] bias_reg_65 = 32'b00000000000000000000000000101011;
reg [32-1:0] bias_reg_66 = 32'b00000000000000000000000001100010;
reg [32-1:0] bias_reg_67 = 32'b00000000000000000000000000010100;
reg [32-1:0] bias_reg_68 = 32'b11111111111111111111111110101110;
reg [32-1:0] bias_reg_69 = 32'b00000000000000000000000000111100;
reg [32-1:0] bias_reg_70 = 32'b11111111111111111111111110011100;
reg [32-1:0] bias_reg_71 = 32'b00000000000000000000000000000111;
reg [32-1:0] bias_reg_72 = 32'b11111111111111111111111111001100;
reg [32-1:0] bias_reg_73 = 32'b11111111111111111111111111010101;
reg [32-1:0] bias_reg_74 = 32'b11111111111111111111111111010000;
reg [32-1:0] bias_reg_75 = 32'b00000000000000000000000010000101;
reg [32-1:0] bias_reg_76 = 32'b11111111111111111111111111011001;
reg [32-1:0] bias_reg_77 = 32'b11111111111111111111111111010101;
reg [32-1:0] bias_reg_78 = 32'b00000000000000000000000000011101;
reg [32-1:0] bias_reg_79 = 32'b11111111111111111111111110011111;
reg [32-1:0] bias_reg_80 = 32'b11111111111111111111111110111110;
reg [32-1:0] bias_reg_81 = 32'b00000000000000000000000000000101;
reg [32-1:0] bias_reg_82 = 32'b11111111111111111111111111100001;
reg [32-1:0] bias_reg_83 = 32'b11111111111111111111111110110000;
reg [32-1:0] bias_reg_84 = 32'b11111111111111111111111111111001;
reg [32-1:0] bias_reg_85 = 32'b11111111111111111111111101111001;
reg [32-1:0] bias_reg_86 = 32'b00000000000000000000000000000011;
reg [32-1:0] bias_reg_87 = 32'b00000000000000000000000100000010;
reg [32-1:0] bias_reg_88 = 32'b11111111111111111111111111101001;
reg [32-1:0] bias_reg_89 = 32'b11111111111111111111111111011101;
reg [32-1:0] bias_reg_90 = 32'b00000000000000000000000001100100;
reg [32-1:0] bias_reg_91 = 32'b11111111111111111111111111000100;
reg [32-1:0] bias_reg_92 = 32'b00000000000000000000000001100001;
reg [32-1:0] bias_reg_93 = 32'b11111111111111111111111110000110;
reg [32-1:0] bias_reg_94 = 32'b11111111111111111111111111000111;
reg [32-1:0] bias_reg_95 = 32'b00000000000000000000000001110001;
reg [32-1:0] bias_reg_96 = 32'b11111111111111111111111111111100;
reg [32-1:0] bias_reg_97 = 32'b00000000000000000000000000110001;
reg [32-1:0] bias_reg_98 = 32'b00000000000000000000000000010101;
reg [32-1:0] bias_reg_99 = 32'b11111111111111111111111111110111;
reg [32-1:0] bias_reg_100 = 32'b00000000000000000000000000000111;
reg [32-1:0] bias_reg_101 = 32'b00000000000000000000000000011000;
reg [32-1:0] bias_reg_102 = 32'b00000000000000000000000000000001;
reg [32-1:0] bias_reg_103 = 32'b11111111111111111111111111000011;
reg [32-1:0] bias_reg_104 = 32'b11111111111111111111111111011111;
reg [32-1:0] bias_reg_105 = 32'b00000000000000000000000010101011;
reg [32-1:0] bias_reg_106 = 32'b00000000000000000000000000110100;
reg [32-1:0] bias_reg_107 = 32'b11111111111111111111111111000111;
reg [32-1:0] bias_reg_108 = 32'b11111111111111111111111111101100;
reg [32-1:0] bias_reg_109 = 32'b11111111111111111111111111110110;
reg [32-1:0] bias_reg_110 = 32'b00000000000000000000000000101111;
reg [32-1:0] bias_reg_111 = 32'b00000000000000000000000001011100;
reg [32-1:0] bias_reg_112 = 32'b00000000000000000000000001011111;
reg [32-1:0] bias_reg_113 = 32'b11111111111111111111111111101111;
reg [32-1:0] bias_reg_114 = 32'b00000000000000000000000001011101;
reg [32-1:0] bias_reg_115 = 32'b11111111111111111111111111110011;
reg [32-1:0] bias_reg_116 = 32'b00000000000000000000000010000011;
reg [32-1:0] bias_reg_117 = 32'b11111111111111111111111111000110;
reg [32-1:0] bias_reg_118 = 32'b00000000000000000000000001000001;
reg [32-1:0] bias_reg_119 = 32'b00000000000000000000000000011001;
reg [32-1:0] bias_reg_120 = 32'b00000000000000000000000000000001;
reg [32-1:0] bias_reg_121 = 32'b11111111111111111111111111001010;
reg [32-1:0] bias_reg_122 = 32'b00000000000000000000000001100001;
reg [32-1:0] bias_reg_123 = 32'b00000000000000000000000001000110;
reg [32-1:0] bias_reg_124 = 32'b00000000000000000000000000100101;
reg [32-1:0] bias_reg_125 = 32'b00000000000000000000000000010100;
reg [32-1:0] bias_reg_126 = 32'b00000000000000000000000001000001;
reg [32-1:0] bias_reg_127 = 32'b11111111111111111111111111101001;
assign bias_mem[0] = bias_reg_0;
assign bias_mem[1] = bias_reg_1;
assign bias_mem[2] = bias_reg_2;
assign bias_mem[3] = bias_reg_3;
assign bias_mem[4] = bias_reg_4;
assign bias_mem[5] = bias_reg_5;
assign bias_mem[6] = bias_reg_6;
assign bias_mem[7] = bias_reg_7;
assign bias_mem[8] = bias_reg_8;
assign bias_mem[9] = bias_reg_9;
assign bias_mem[10] = bias_reg_10;
assign bias_mem[11] = bias_reg_11;
assign bias_mem[12] = bias_reg_12;
assign bias_mem[13] = bias_reg_13;
assign bias_mem[14] = bias_reg_14;
assign bias_mem[15] = bias_reg_15;
assign bias_mem[16] = bias_reg_16;
assign bias_mem[17] = bias_reg_17;
assign bias_mem[18] = bias_reg_18;
assign bias_mem[19] = bias_reg_19;
assign bias_mem[20] = bias_reg_20;
assign bias_mem[21] = bias_reg_21;
assign bias_mem[22] = bias_reg_22;
assign bias_mem[23] = bias_reg_23;
assign bias_mem[24] = bias_reg_24;
assign bias_mem[25] = bias_reg_25;
assign bias_mem[26] = bias_reg_26;
assign bias_mem[27] = bias_reg_27;
assign bias_mem[28] = bias_reg_28;
assign bias_mem[29] = bias_reg_29;
assign bias_mem[30] = bias_reg_30;
assign bias_mem[31] = bias_reg_31;
assign bias_mem[32] = bias_reg_32;
assign bias_mem[33] = bias_reg_33;
assign bias_mem[34] = bias_reg_34;
assign bias_mem[35] = bias_reg_35;
assign bias_mem[36] = bias_reg_36;
assign bias_mem[37] = bias_reg_37;
assign bias_mem[38] = bias_reg_38;
assign bias_mem[39] = bias_reg_39;
assign bias_mem[40] = bias_reg_40;
assign bias_mem[41] = bias_reg_41;
assign bias_mem[42] = bias_reg_42;
assign bias_mem[43] = bias_reg_43;
assign bias_mem[44] = bias_reg_44;
assign bias_mem[45] = bias_reg_45;
assign bias_mem[46] = bias_reg_46;
assign bias_mem[47] = bias_reg_47;
assign bias_mem[48] = bias_reg_48;
assign bias_mem[49] = bias_reg_49;
assign bias_mem[50] = bias_reg_50;
assign bias_mem[51] = bias_reg_51;
assign bias_mem[52] = bias_reg_52;
assign bias_mem[53] = bias_reg_53;
assign bias_mem[54] = bias_reg_54;
assign bias_mem[55] = bias_reg_55;
assign bias_mem[56] = bias_reg_56;
assign bias_mem[57] = bias_reg_57;
assign bias_mem[58] = bias_reg_58;
assign bias_mem[59] = bias_reg_59;
assign bias_mem[60] = bias_reg_60;
assign bias_mem[61] = bias_reg_61;
assign bias_mem[62] = bias_reg_62;
assign bias_mem[63] = bias_reg_63;
assign bias_mem[64] = bias_reg_64;
assign bias_mem[65] = bias_reg_65;
assign bias_mem[66] = bias_reg_66;
assign bias_mem[67] = bias_reg_67;
assign bias_mem[68] = bias_reg_68;
assign bias_mem[69] = bias_reg_69;
assign bias_mem[70] = bias_reg_70;
assign bias_mem[71] = bias_reg_71;
assign bias_mem[72] = bias_reg_72;
assign bias_mem[73] = bias_reg_73;
assign bias_mem[74] = bias_reg_74;
assign bias_mem[75] = bias_reg_75;
assign bias_mem[76] = bias_reg_76;
assign bias_mem[77] = bias_reg_77;
assign bias_mem[78] = bias_reg_78;
assign bias_mem[79] = bias_reg_79;
assign bias_mem[80] = bias_reg_80;
assign bias_mem[81] = bias_reg_81;
assign bias_mem[82] = bias_reg_82;
assign bias_mem[83] = bias_reg_83;
assign bias_mem[84] = bias_reg_84;
assign bias_mem[85] = bias_reg_85;
assign bias_mem[86] = bias_reg_86;
assign bias_mem[87] = bias_reg_87;
assign bias_mem[88] = bias_reg_88;
assign bias_mem[89] = bias_reg_89;
assign bias_mem[90] = bias_reg_90;
assign bias_mem[91] = bias_reg_91;
assign bias_mem[92] = bias_reg_92;
assign bias_mem[93] = bias_reg_93;
assign bias_mem[94] = bias_reg_94;
assign bias_mem[95] = bias_reg_95;
assign bias_mem[96] = bias_reg_96;
assign bias_mem[97] = bias_reg_97;
assign bias_mem[98] = bias_reg_98;
assign bias_mem[99] = bias_reg_99;
assign bias_mem[100] = bias_reg_100;
assign bias_mem[101] = bias_reg_101;
assign bias_mem[102] = bias_reg_102;
assign bias_mem[103] = bias_reg_103;
assign bias_mem[104] = bias_reg_104;
assign bias_mem[105] = bias_reg_105;
assign bias_mem[106] = bias_reg_106;
assign bias_mem[107] = bias_reg_107;
assign bias_mem[108] = bias_reg_108;
assign bias_mem[109] = bias_reg_109;
assign bias_mem[110] = bias_reg_110;
assign bias_mem[111] = bias_reg_111;
assign bias_mem[112] = bias_reg_112;
assign bias_mem[113] = bias_reg_113;
assign bias_mem[114] = bias_reg_114;
assign bias_mem[115] = bias_reg_115;
assign bias_mem[116] = bias_reg_116;
assign bias_mem[117] = bias_reg_117;
assign bias_mem[118] = bias_reg_118;
assign bias_mem[119] = bias_reg_119;
assign bias_mem[120] = bias_reg_120;
assign bias_mem[121] = bias_reg_121;
assign bias_mem[122] = bias_reg_122;
assign bias_mem[123] = bias_reg_123;
assign bias_mem[124] = bias_reg_124;
assign bias_mem[125] = bias_reg_125;
assign bias_mem[126] = bias_reg_126;
assign bias_mem[127] = bias_reg_127;
endmodule
