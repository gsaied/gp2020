/*
* FIRE2 SQUEEZE 3*3 IMPLEMENTATION
* INPUT SIZE: 128*128*64
* OUTPUT SIZE: 64*64*16
* STRIDE: 1
* PAD:	1
* WINDOW: 3*3
*/
module fire2_squeeze_3 #(
	parameter WOUT = 64 ,
	parameter DSP_NO = 16,
	parameter STRIDE = 2 ,
	parameter W_IN = 128,
	parameter WIDTH = 16 ,
	parameter CHIN = 64 , 
	parameter KERNEL_DIM = 3 ,
	parameter CHOUT = 16   
)
(
	input clk,
	input rst,
	input fire2_squeeze_3_en,
	output reg fire2_squeeze_3_sample,
	input [15:0] ifm,
	output reg fire2_squeeze_3_end,
	output reg [WIDTH-1:0] ofm [0:DSP_NO-1]
);

wire [2*WIDTH-1:0] biasing_wire [0:DSP_NO-1] ;
biasing_rom b7 (
	.bias_mem(biasing_wire)
);
///////////////////////////////////
//KERNELS INSTANTIATION
///////////////////////////////////
wire [WIDTH-1:0] kernels [0:DSP_NO-1] ; 
//reg [WIDTH-1:0] kernel_regs [0:DSP_NO-1] ; 
reg [$clog2(CHIN*KERNEL_DIM**2)-1:0] weight_rom_address ; 
//////////////////////////////////
rom_array_layer_1 u_2 (
	.clk(clk),
	.address(weight_rom_address),
	.rom_out(kernels)
);
///////////////////////////////////
//this signal is very important to track
//represents a pulse to clr pin of mac to reset every 27 cycles of clk
///////////////////////////////////
reg clr_pulse ; 
///////
///////
always @(posedge clk or negedge rst) begin
	if(!rst)
		weight_rom_address<= 0 ; 
	else if (rom_clr_pulse)
		weight_rom_address<= 0;
	else begin
		weight_rom_address<= weight_rom_address+1;
	end
end
reg rom_clr_pulse ; 
/*
always @(posedge clk) begin
	kernel_regs<=kernels ;		
end
*/
////////////////////////////
//GENERATION OF CLR PULSE///
////////////////////////////
reg [$clog2(KERNEL_DIM**2*CHIN):0] counter_10 ; 
always @(posedge clk or negedge rst) begin
	if(!rst) begin
		clr_pulse <= 1'b0 ; 
		rom_clr_pulse <= 1'b0 ; 
		counter_10 <= 0 ;
	end
	else if (!fire2_squeeze_3_end) begin
		if(counter_10 == KERNEL_DIM**2*CHIN) begin
			counter_10 <= 0 ;
			clr_pulse<= 1'b1 ;
			rom_clr_pulse<= 1'b0 ; 
		end
		else if(counter_10 == KERNEL_DIM**2*CHIN-1) begin
			counter_10 <= counter_10+1  ;
			rom_clr_pulse<= 1'b1 ;
		end
		else begin
			clr_pulse <= 1'b0 ; 
			rom_clr_pulse<= 1'b0 ; 
			counter_10 <= counter_10 +1;
		end
	end
end
//////////////////////////////
//CORE GENERATION/////////////
//////////////////////////////
wire [2*WIDTH:0] ofmw [0:DSP_NO-1];
reg [2*WIDTH:0] ofmw2 [0:DSP_NO-1];
genvar i ; 
generate for (i = 0 ; i< CHOUT ; i++) begin
	mac mac_i (
		.clr(clr_pulse),
		.clk(clk),
		.rst(rst),
		.pix(ifm),
		.mul_out(ofmw[i]),
		.ker(kernels[i])
	);
end
endgenerate
/////////////////////////////////
//OUTPUT IS READY TO BE SAMPLED//
/////////////////////////////////
always @(*) begin
	for (int i = 0 ; i < DSP_NO ; i++) begin
		ofmw2[i]  = ofmw[i] + biasing_wire[i]  ;
	end
end
always@(posedge clk) begin
	if(fire2_squeeze_3_en && !fire2_squeeze_3_end && clr_pulse) begin
		for (int i = 0 ; i< DSP_NO ; i++) begin
			if(ofmw2[i][31] == 1'b1 || ofmw2[i][32] == 1'b1 ) 
				ofm[i] <= 16'b0 ;
			else
				ofm[i] <= {ofmw2[i][31],ofmw2[i][28:14]};
		end
	end
end
///////////////////////////////
//CHECK FOR LAYER END//////////
///////////////////////////////
reg [$clog2(WOUT**2):0] fire2_squeeze_3_timer ;// will be changed
always @(posedge clk or negedge rst) begin
	if (!rst) begin
		fire2_squeeze_3_timer<= 0 ;
		fire2_squeeze_3_end <= 1'b0 ; 
	end
	else if (fire2_squeeze_3_timer == WOUT**2)// will be changed
		fire2_squeeze_3_end <= 1'b1 ;//LAYER_1 HAS FINISHED
	else if (clr_pulse)
		fire2_squeeze_3_timer<= fire2_squeeze_3_timer+1 ; 

end
always @(posedge clk) begin
   fire2_squeeze_3_sample <= clr_pulse ;
end
endmodule

