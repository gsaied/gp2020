
	/* verilator lint_off COMBDLY */
	module rom_3 #(
	parameter WIDTH=16,
	parameter KERNEL=1,
	parameter ADDR=4,
	parameter NUM=64)
	(
		input [ADDR-1:0] address ,
		input clk,
		output reg [WIDTH-1:0] rom_out [0:NUM-1]
	);	
	

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_1 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_2 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_3 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_4 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_5 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_6 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_7 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_8 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_9 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_10 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_11 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_12 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_13 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_14 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_15 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_16 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_17 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_18 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_19 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_20 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_21 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_22 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_23 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_24 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_25 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_26 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_27 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_28 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_29 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_30 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_31 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_32 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_33 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_34 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_35 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_36 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_37 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_38 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_39 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_40 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_41 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_42 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_43 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_44 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_45 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_46 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_47 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_48 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_49 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_50 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_51 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_52 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_53 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_54 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_55 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_56 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_57 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_58 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_59 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_60 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_61 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_62 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_63 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_64 [0:2**ADDR-1] ;
initial  begin
$readmemb("file_1_2.mem",rom_1,0,16-1);
$readmemb("file_2_2.mem",rom_2,0,2**ADDR-1);
$readmemb("file_3_2.mem",rom_3,0,2**ADDR-1);
$readmemb("file_4_2.mem",rom_4,0,2**ADDR-1);
$readmemb("file_5_2.mem",rom_5,0,2**ADDR-1);
$readmemb("file_6_2.mem",rom_6,0,2**ADDR-1);
$readmemb("file_7_2.mem",rom_7,0,2**ADDR-1);
$readmemb("file_8_2.mem",rom_8,0,2**ADDR-1);
$readmemb("file_9_2.mem",rom_9,0,2**ADDR-1);
$readmemb("file_10_2.mem",rom_10,0,2**ADDR-1);
$readmemb("file_11_2.mem",rom_11,0,2**ADDR-1);
$readmemb("file_12_2.mem",rom_12,0,2**ADDR-1);
$readmemb("file_13_2.mem",rom_13,0,2**ADDR-1);
$readmemb("file_14_2.mem",rom_14,0,2**ADDR-1);
$readmemb("file_15_2.mem",rom_15,0,2**ADDR-1);
$readmemb("file_16_2.mem",rom_16,0,2**ADDR-1);
$readmemb("file_17_2.mem",rom_17,0,2**ADDR-1);
$readmemb("file_18_2.mem",rom_18,0,2**ADDR-1);
$readmemb("file_19_2.mem",rom_19,0,2**ADDR-1);
$readmemb("file_20_2.mem",rom_20,0,2**ADDR-1);
$readmemb("file_21_2.mem",rom_21,0,2**ADDR-1);
$readmemb("file_22_2.mem",rom_22,0,2**ADDR-1);
$readmemb("file_23_2.mem",rom_23,0,2**ADDR-1);
$readmemb("file_24_2.mem",rom_24,0,2**ADDR-1);
$readmemb("file_25_2.mem",rom_25,0,2**ADDR-1);
$readmemb("file_26_2.mem",rom_26,0,2**ADDR-1);
$readmemb("file_27_2.mem",rom_27,0,2**ADDR-1);
$readmemb("file_28_2.mem",rom_28,0,2**ADDR-1);
$readmemb("file_29_2.mem",rom_29,0,2**ADDR-1);
$readmemb("file_30_2.mem",rom_30,0,2**ADDR-1);
$readmemb("file_31_2.mem",rom_31,0,2**ADDR-1);
$readmemb("file_32_2.mem",rom_32,0,2**ADDR-1);
$readmemb("file_33_2.mem",rom_33,0,2**ADDR-1);
$readmemb("file_34_2.mem",rom_34,0,2**ADDR-1);
$readmemb("file_35_2.mem",rom_35,0,2**ADDR-1);
$readmemb("file_36_2.mem",rom_36,0,2**ADDR-1);
$readmemb("file_37_2.mem",rom_37,0,2**ADDR-1);
$readmemb("file_38_2.mem",rom_38,0,2**ADDR-1);
$readmemb("file_39_2.mem",rom_39,0,2**ADDR-1);
$readmemb("file_40_2.mem",rom_40,0,2**ADDR-1);
$readmemb("file_41_2.mem",rom_41,0,2**ADDR-1);
$readmemb("file_42_2.mem",rom_42,0,2**ADDR-1);
$readmemb("file_43_2.mem",rom_43,0,2**ADDR-1);
$readmemb("file_44_2.mem",rom_44,0,2**ADDR-1);
$readmemb("file_45_2.mem",rom_45,0,2**ADDR-1);
$readmemb("file_46_2.mem",rom_46,0,2**ADDR-1);
$readmemb("file_47_2.mem",rom_47,0,2**ADDR-1);
$readmemb("file_48_2.mem",rom_48,0,2**ADDR-1);
$readmemb("file_49_2.mem",rom_49,0,2**ADDR-1);
$readmemb("file_50_2.mem",rom_50,0,2**ADDR-1);
$readmemb("file_51_2.mem",rom_51,0,2**ADDR-1);
$readmemb("file_52_2.mem",rom_52,0,2**ADDR-1);
$readmemb("file_53_2.mem",rom_53,0,2**ADDR-1);
$readmemb("file_54_2.mem",rom_54,0,2**ADDR-1);
$readmemb("file_55_2.mem",rom_55,0,2**ADDR-1);
$readmemb("file_56_2.mem",rom_56,0,2**ADDR-1);
$readmemb("file_57_2.mem",rom_57,0,2**ADDR-1);
$readmemb("file_58_2.mem",rom_58,0,2**ADDR-1);
$readmemb("file_59_2.mem",rom_59,0,2**ADDR-1);
$readmemb("file_60_2.mem",rom_60,0,2**ADDR-1);
$readmemb("file_61_2.mem",rom_61,0,2**ADDR-1);
$readmemb("file_62_2.mem",rom_62,0,2**ADDR-1);
$readmemb("file_63_2.mem",rom_63,0,2**ADDR-1);
$readmemb("file_64_2.mem",rom_64,0,2**ADDR-1);
end
always @(posedge clk ) begin
 rom_out[0]<= rom_1[address] ;
 rom_out[1]<= rom_2[address] ;
 rom_out[2]<= rom_3[address] ;
 rom_out[3]<= rom_4[address] ;
 rom_out[4]<= rom_5[address] ;
 rom_out[5]<= rom_6[address] ;
 rom_out[6]<= rom_7[address] ;
 rom_out[7]<= rom_8[address] ;
 rom_out[8]<= rom_9[address] ;
 rom_out[9]<= rom_10[address] ;
 rom_out[10]<= rom_11[address] ;
 rom_out[11]<= rom_12[address] ;
 rom_out[12]<= rom_13[address] ;
 rom_out[13]<= rom_14[address] ;
 rom_out[14]<= rom_15[address] ;
 rom_out[15]<= rom_16[address] ;
 rom_out[16]<= rom_17[address] ;
 rom_out[17]<= rom_18[address] ;
 rom_out[18]<= rom_19[address] ;
 rom_out[19]<= rom_20[address] ;
 rom_out[20]<= rom_21[address] ;
 rom_out[21]<= rom_22[address] ;
 rom_out[22]<= rom_23[address] ;
 rom_out[23]<= rom_24[address] ;
 rom_out[24]<= rom_25[address] ;
 rom_out[25]<= rom_26[address] ;
 rom_out[26]<= rom_27[address] ;
 rom_out[27]<= rom_28[address] ;
 rom_out[28]<= rom_29[address] ;
 rom_out[29]<= rom_30[address] ;
 rom_out[30]<= rom_31[address] ;
 rom_out[31]<= rom_32[address] ;
 rom_out[32]<= rom_33[address] ;
 rom_out[33]<= rom_34[address] ;
 rom_out[34]<= rom_35[address] ;
 rom_out[35]<= rom_36[address] ;
 rom_out[36]<= rom_37[address] ;
 rom_out[37]<= rom_38[address] ;
 rom_out[38]<= rom_39[address] ;
 rom_out[39]<= rom_40[address] ;
 rom_out[40]<= rom_41[address] ;
 rom_out[41]<= rom_42[address] ;
 rom_out[42]<= rom_43[address] ;
 rom_out[43]<= rom_44[address] ;
 rom_out[44]<= rom_45[address] ;
 rom_out[45]<= rom_46[address] ;
 rom_out[46]<= rom_47[address] ;
 rom_out[47]<= rom_48[address] ;
 rom_out[48]<= rom_49[address] ;
 rom_out[49]<= rom_50[address] ;
 rom_out[50]<= rom_51[address] ;
 rom_out[51]<= rom_52[address] ;
 rom_out[52]<= rom_53[address] ;
 rom_out[53]<= rom_54[address] ;
 rom_out[54]<= rom_55[address] ;
 rom_out[55]<= rom_56[address] ;
 rom_out[56]<= rom_57[address] ;
 rom_out[57]<= rom_58[address] ;
 rom_out[58]<= rom_59[address] ;
 rom_out[59]<= rom_60[address] ;
 rom_out[60]<= rom_61[address] ;
 rom_out[61]<= rom_62[address] ;
 rom_out[62]<= rom_63[address] ;
 rom_out[63]<= rom_64[address] ;
end
endmodule
